module alu_4 (A,
    B,
    CTRL,
    Y);
 input [3:0] A;
 input [3:0] B;
 input [3:0] CTRL;
 output [7:0] Y;

 wire VDD;
 wire VSS;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _130_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_127 ();
 FILLCELL_X32 FILLER_0_159 ();
 FILLCELL_X8 FILLER_0_17 ();
 FILLCELL_X32 FILLER_0_191 ();
 FILLCELL_X16 FILLER_0_223 ();
 FILLCELL_X4 FILLER_0_239 ();
 FILLCELL_X1 FILLER_0_243 ();
 FILLCELL_X1 FILLER_0_244 ();
 FILLCELL_X1 FILLER_0_29 ();
 FILLCELL_X1 FILLER_0_30 ();
 FILLCELL_X16 FILLER_0_34 ();
 FILLCELL_X1 FILLER_0_50 ();
 FILLCELL_X1 FILLER_0_51 ();
 FILLCELL_X1 FILLER_0_52 ();
 FILLCELL_X1 FILLER_0_57 ();
 FILLCELL_X1 FILLER_0_58 ();
 FILLCELL_X32 FILLER_0_63 ();
 FILLCELL_X32 FILLER_0_95 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X4 FILLER_10_111 ();
 FILLCELL_X4 FILLER_10_118 ();
 FILLCELL_X1 FILLER_10_122 ();
 FILLCELL_X32 FILLER_10_125 ();
 FILLCELL_X32 FILLER_10_157 ();
 FILLCELL_X8 FILLER_10_17 ();
 FILLCELL_X32 FILLER_10_189 ();
 FILLCELL_X16 FILLER_10_221 ();
 FILLCELL_X8 FILLER_10_237 ();
 FILLCELL_X4 FILLER_10_25 ();
 FILLCELL_X1 FILLER_10_29 ();
 FILLCELL_X1 FILLER_10_30 ();
 FILLCELL_X8 FILLER_10_41 ();
 FILLCELL_X4 FILLER_10_49 ();
 FILLCELL_X1 FILLER_10_53 ();
 FILLCELL_X1 FILLER_10_54 ();
 FILLCELL_X8 FILLER_10_58 ();
 FILLCELL_X4 FILLER_10_66 ();
 FILLCELL_X1 FILLER_10_72 ();
 FILLCELL_X1 FILLER_10_73 ();
 FILLCELL_X4 FILLER_10_78 ();
 FILLCELL_X4 FILLER_10_85 ();
 FILLCELL_X1 FILLER_10_89 ();
 FILLCELL_X1 FILLER_10_90 ();
 FILLCELL_X16 FILLER_10_95 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X1 FILLER_11_102 ();
 FILLCELL_X16 FILLER_11_106 ();
 FILLCELL_X8 FILLER_11_122 ();
 FILLCELL_X4 FILLER_11_130 ();
 FILLCELL_X32 FILLER_11_137 ();
 FILLCELL_X8 FILLER_11_169 ();
 FILLCELL_X4 FILLER_11_177 ();
 FILLCELL_X1 FILLER_11_181 ();
 FILLCELL_X1 FILLER_11_182 ();
 FILLCELL_X1 FILLER_11_186 ();
 FILLCELL_X1 FILLER_11_187 ();
 FILLCELL_X8 FILLER_11_191 ();
 FILLCELL_X1 FILLER_11_199 ();
 FILLCELL_X1 FILLER_11_200 ();
 FILLCELL_X1 FILLER_11_217 ();
 FILLCELL_X1 FILLER_11_218 ();
 FILLCELL_X1 FILLER_11_222 ();
 FILLCELL_X1 FILLER_11_223 ();
 FILLCELL_X8 FILLER_11_227 ();
 FILLCELL_X4 FILLER_11_235 ();
 FILLCELL_X1 FILLER_11_239 ();
 FILLCELL_X1 FILLER_11_243 ();
 FILLCELL_X1 FILLER_11_244 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X4 FILLER_11_65 ();
 FILLCELL_X1 FILLER_11_69 ();
 FILLCELL_X1 FILLER_11_70 ();
 FILLCELL_X16 FILLER_11_74 ();
 FILLCELL_X8 FILLER_11_90 ();
 FILLCELL_X4 FILLER_11_98 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X16 FILLER_12_115 ();
 FILLCELL_X4 FILLER_12_131 ();
 FILLCELL_X1 FILLER_12_135 ();
 FILLCELL_X1 FILLER_12_139 ();
 FILLCELL_X1 FILLER_12_140 ();
 FILLCELL_X16 FILLER_12_144 ();
 FILLCELL_X8 FILLER_12_160 ();
 FILLCELL_X4 FILLER_12_17 ();
 FILLCELL_X16 FILLER_12_184 ();
 FILLCELL_X8 FILLER_12_200 ();
 FILLCELL_X1 FILLER_12_208 ();
 FILLCELL_X1 FILLER_12_209 ();
 FILLCELL_X1 FILLER_12_214 ();
 FILLCELL_X1 FILLER_12_215 ();
 FILLCELL_X16 FILLER_12_220 ();
 FILLCELL_X4 FILLER_12_23 ();
 FILLCELL_X8 FILLER_12_236 ();
 FILLCELL_X1 FILLER_12_244 ();
 FILLCELL_X16 FILLER_12_29 ();
 FILLCELL_X8 FILLER_12_45 ();
 FILLCELL_X4 FILLER_12_53 ();
 FILLCELL_X16 FILLER_12_60 ();
 FILLCELL_X1 FILLER_12_76 ();
 FILLCELL_X1 FILLER_12_77 ();
 FILLCELL_X1 FILLER_12_78 ();
 FILLCELL_X32 FILLER_12_83 ();
 FILLCELL_X16 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_103 ();
 FILLCELL_X8 FILLER_13_135 ();
 FILLCELL_X4 FILLER_13_143 ();
 FILLCELL_X1 FILLER_13_147 ();
 FILLCELL_X1 FILLER_13_148 ();
 FILLCELL_X16 FILLER_13_153 ();
 FILLCELL_X4 FILLER_13_169 ();
 FILLCELL_X8 FILLER_13_17 ();
 FILLCELL_X1 FILLER_13_173 ();
 FILLCELL_X32 FILLER_13_177 ();
 FILLCELL_X8 FILLER_13_209 ();
 FILLCELL_X1 FILLER_13_217 ();
 FILLCELL_X1 FILLER_13_218 ();
 FILLCELL_X16 FILLER_13_222 ();
 FILLCELL_X1 FILLER_13_238 ();
 FILLCELL_X1 FILLER_13_239 ();
 FILLCELL_X1 FILLER_13_243 ();
 FILLCELL_X1 FILLER_13_244 ();
 FILLCELL_X1 FILLER_13_25 ();
 FILLCELL_X1 FILLER_13_26 ();
 FILLCELL_X1 FILLER_13_27 ();
 FILLCELL_X1 FILLER_13_30 ();
 FILLCELL_X1 FILLER_13_31 ();
 FILLCELL_X8 FILLER_13_34 ();
 FILLCELL_X4 FILLER_13_42 ();
 FILLCELL_X1 FILLER_13_46 ();
 FILLCELL_X1 FILLER_13_47 ();
 FILLCELL_X1 FILLER_13_48 ();
 FILLCELL_X4 FILLER_13_53 ();
 FILLCELL_X16 FILLER_13_61 ();
 FILLCELL_X8 FILLER_13_77 ();
 FILLCELL_X4 FILLER_13_85 ();
 FILLCELL_X1 FILLER_13_89 ();
 FILLCELL_X1 FILLER_13_92 ();
 FILLCELL_X1 FILLER_13_93 ();
 FILLCELL_X4 FILLER_13_97 ();
 FILLCELL_X8 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_100 ();
 FILLCELL_X16 FILLER_14_103 ();
 FILLCELL_X8 FILLER_14_119 ();
 FILLCELL_X4 FILLER_14_127 ();
 FILLCELL_X1 FILLER_14_13 ();
 FILLCELL_X1 FILLER_14_131 ();
 FILLCELL_X1 FILLER_14_132 ();
 FILLCELL_X1 FILLER_14_133 ();
 FILLCELL_X8 FILLER_14_136 ();
 FILLCELL_X1 FILLER_14_14 ();
 FILLCELL_X1 FILLER_14_144 ();
 FILLCELL_X1 FILLER_14_149 ();
 FILLCELL_X1 FILLER_14_150 ();
 FILLCELL_X4 FILLER_14_161 ();
 FILLCELL_X1 FILLER_14_165 ();
 FILLCELL_X1 FILLER_14_169 ();
 FILLCELL_X1 FILLER_14_170 ();
 FILLCELL_X1 FILLER_14_171 ();
 FILLCELL_X8 FILLER_14_175 ();
 FILLCELL_X1 FILLER_14_183 ();
 FILLCELL_X1 FILLER_14_184 ();
 FILLCELL_X16 FILLER_14_187 ();
 FILLCELL_X4 FILLER_14_203 ();
 FILLCELL_X1 FILLER_14_207 ();
 FILLCELL_X1 FILLER_14_208 ();
 FILLCELL_X1 FILLER_14_212 ();
 FILLCELL_X1 FILLER_14_213 ();
 FILLCELL_X1 FILLER_14_217 ();
 FILLCELL_X1 FILLER_14_218 ();
 FILLCELL_X16 FILLER_14_222 ();
 FILLCELL_X4 FILLER_14_238 ();
 FILLCELL_X1 FILLER_14_242 ();
 FILLCELL_X1 FILLER_14_243 ();
 FILLCELL_X1 FILLER_14_244 ();
 FILLCELL_X1 FILLER_14_25 ();
 FILLCELL_X1 FILLER_14_26 ();
 FILLCELL_X32 FILLER_14_43 ();
 FILLCELL_X1 FILLER_14_75 ();
 FILLCELL_X4 FILLER_14_9 ();
 FILLCELL_X8 FILLER_14_92 ();
 FILLCELL_X16 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_100 ();
 FILLCELL_X1 FILLER_15_101 ();
 FILLCELL_X1 FILLER_15_105 ();
 FILLCELL_X1 FILLER_15_106 ();
 FILLCELL_X32 FILLER_15_110 ();
 FILLCELL_X4 FILLER_15_142 ();
 FILLCELL_X1 FILLER_15_146 ();
 FILLCELL_X32 FILLER_15_163 ();
 FILLCELL_X4 FILLER_15_17 ();
 FILLCELL_X1 FILLER_15_195 ();
 FILLCELL_X1 FILLER_15_196 ();
 FILLCELL_X1 FILLER_15_197 ();
 FILLCELL_X1 FILLER_15_200 ();
 FILLCELL_X1 FILLER_15_201 ();
 FILLCELL_X16 FILLER_15_218 ();
 FILLCELL_X8 FILLER_15_23 ();
 FILLCELL_X8 FILLER_15_234 ();
 FILLCELL_X1 FILLER_15_242 ();
 FILLCELL_X1 FILLER_15_243 ();
 FILLCELL_X1 FILLER_15_244 ();
 FILLCELL_X1 FILLER_15_31 ();
 FILLCELL_X32 FILLER_15_42 ();
 FILLCELL_X16 FILLER_15_74 ();
 FILLCELL_X1 FILLER_15_90 ();
 FILLCELL_X1 FILLER_15_91 ();
 FILLCELL_X1 FILLER_15_92 ();
 FILLCELL_X4 FILLER_15_96 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_100 ();
 FILLCELL_X16 FILLER_16_132 ();
 FILLCELL_X1 FILLER_16_158 ();
 FILLCELL_X1 FILLER_16_159 ();
 FILLCELL_X32 FILLER_16_162 ();
 FILLCELL_X8 FILLER_16_194 ();
 FILLCELL_X1 FILLER_16_202 ();
 FILLCELL_X1 FILLER_16_203 ();
 FILLCELL_X1 FILLER_16_204 ();
 FILLCELL_X32 FILLER_16_208 ();
 FILLCELL_X4 FILLER_16_240 ();
 FILLCELL_X1 FILLER_16_244 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X16 FILLER_16_65 ();
 FILLCELL_X4 FILLER_16_81 ();
 FILLCELL_X1 FILLER_16_85 ();
 FILLCELL_X1 FILLER_16_96 ();
 FILLCELL_X1 FILLER_16_97 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_123 ();
 FILLCELL_X32 FILLER_17_155 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X16 FILLER_17_187 ();
 FILLCELL_X1 FILLER_17_203 ();
 FILLCELL_X16 FILLER_17_214 ();
 FILLCELL_X8 FILLER_17_230 ();
 FILLCELL_X4 FILLER_17_238 ();
 FILLCELL_X1 FILLER_17_242 ();
 FILLCELL_X1 FILLER_17_243 ();
 FILLCELL_X1 FILLER_17_244 ();
 FILLCELL_X32 FILLER_17_27 ();
 FILLCELL_X32 FILLER_17_59 ();
 FILLCELL_X32 FILLER_17_91 ();
 FILLCELL_X8 FILLER_18_1 ();
 FILLCELL_X4 FILLER_18_121 ();
 FILLCELL_X1 FILLER_18_125 ();
 FILLCELL_X1 FILLER_18_126 ();
 FILLCELL_X1 FILLER_18_127 ();
 FILLCELL_X1 FILLER_18_13 ();
 FILLCELL_X16 FILLER_18_130 ();
 FILLCELL_X1 FILLER_18_14 ();
 FILLCELL_X8 FILLER_18_146 ();
 FILLCELL_X4 FILLER_18_154 ();
 FILLCELL_X1 FILLER_18_158 ();
 FILLCELL_X1 FILLER_18_159 ();
 FILLCELL_X1 FILLER_18_160 ();
 FILLCELL_X32 FILLER_18_164 ();
 FILLCELL_X1 FILLER_18_18 ();
 FILLCELL_X1 FILLER_18_19 ();
 FILLCELL_X8 FILLER_18_196 ();
 FILLCELL_X4 FILLER_18_204 ();
 FILLCELL_X16 FILLER_18_224 ();
 FILLCELL_X1 FILLER_18_23 ();
 FILLCELL_X1 FILLER_18_24 ();
 FILLCELL_X4 FILLER_18_240 ();
 FILLCELL_X1 FILLER_18_244 ();
 FILLCELL_X1 FILLER_18_27 ();
 FILLCELL_X1 FILLER_18_28 ();
 FILLCELL_X32 FILLER_18_39 ();
 FILLCELL_X16 FILLER_18_71 ();
 FILLCELL_X32 FILLER_18_89 ();
 FILLCELL_X4 FILLER_18_9 ();
 FILLCELL_X1 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_104 ();
 FILLCELL_X32 FILLER_19_136 ();
 FILLCELL_X32 FILLER_19_168 ();
 FILLCELL_X1 FILLER_19_2 ();
 FILLCELL_X8 FILLER_19_200 ();
 FILLCELL_X1 FILLER_19_208 ();
 FILLCELL_X1 FILLER_19_209 ();
 FILLCELL_X1 FILLER_19_210 ();
 FILLCELL_X32 FILLER_19_213 ();
 FILLCELL_X8 FILLER_19_23 ();
 FILLCELL_X4 FILLER_19_31 ();
 FILLCELL_X1 FILLER_19_35 ();
 FILLCELL_X1 FILLER_19_36 ();
 FILLCELL_X1 FILLER_19_37 ();
 FILLCELL_X32 FILLER_19_40 ();
 FILLCELL_X16 FILLER_19_7 ();
 FILLCELL_X32 FILLER_19_72 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X4 FILLER_1_101 ();
 FILLCELL_X1 FILLER_1_105 ();
 FILLCELL_X1 FILLER_1_106 ();
 FILLCELL_X32 FILLER_1_110 ();
 FILLCELL_X32 FILLER_1_142 ();
 FILLCELL_X8 FILLER_1_17 ();
 FILLCELL_X32 FILLER_1_174 ();
 FILLCELL_X32 FILLER_1_206 ();
 FILLCELL_X1 FILLER_1_238 ();
 FILLCELL_X1 FILLER_1_239 ();
 FILLCELL_X1 FILLER_1_243 ();
 FILLCELL_X1 FILLER_1_244 ();
 FILLCELL_X4 FILLER_1_25 ();
 FILLCELL_X32 FILLER_1_32 ();
 FILLCELL_X32 FILLER_1_64 ();
 FILLCELL_X1 FILLER_1_96 ();
 FILLCELL_X1 FILLER_1_97 ();
 FILLCELL_X1 FILLER_20_1 ();
 FILLCELL_X4 FILLER_20_105 ();
 FILLCELL_X1 FILLER_20_109 ();
 FILLCELL_X1 FILLER_20_110 ();
 FILLCELL_X1 FILLER_20_111 ();
 FILLCELL_X1 FILLER_20_122 ();
 FILLCELL_X1 FILLER_20_123 ();
 FILLCELL_X4 FILLER_20_126 ();
 FILLCELL_X1 FILLER_20_130 ();
 FILLCELL_X1 FILLER_20_131 ();
 FILLCELL_X1 FILLER_20_132 ();
 FILLCELL_X8 FILLER_20_14 ();
 FILLCELL_X8 FILLER_20_149 ();
 FILLCELL_X4 FILLER_20_157 ();
 FILLCELL_X1 FILLER_20_161 ();
 FILLCELL_X1 FILLER_20_162 ();
 FILLCELL_X1 FILLER_20_163 ();
 FILLCELL_X1 FILLER_20_174 ();
 FILLCELL_X1 FILLER_20_175 ();
 FILLCELL_X1 FILLER_20_176 ();
 FILLCELL_X8 FILLER_20_179 ();
 FILLCELL_X4 FILLER_20_187 ();
 FILLCELL_X1 FILLER_20_191 ();
 FILLCELL_X1 FILLER_20_194 ();
 FILLCELL_X1 FILLER_20_195 ();
 FILLCELL_X1 FILLER_20_199 ();
 FILLCELL_X1 FILLER_20_2 ();
 FILLCELL_X1 FILLER_20_200 ();
 FILLCELL_X16 FILLER_20_217 ();
 FILLCELL_X8 FILLER_20_233 ();
 FILLCELL_X4 FILLER_20_241 ();
 FILLCELL_X4 FILLER_20_25 ();
 FILLCELL_X1 FILLER_20_29 ();
 FILLCELL_X1 FILLER_20_30 ();
 FILLCELL_X1 FILLER_20_31 ();
 FILLCELL_X8 FILLER_20_48 ();
 FILLCELL_X1 FILLER_20_56 ();
 FILLCELL_X1 FILLER_20_57 ();
 FILLCELL_X4 FILLER_20_60 ();
 FILLCELL_X1 FILLER_20_64 ();
 FILLCELL_X1 FILLER_20_65 ();
 FILLCELL_X1 FILLER_20_68 ();
 FILLCELL_X1 FILLER_20_69 ();
 FILLCELL_X1 FILLER_20_8 ();
 FILLCELL_X1 FILLER_20_80 ();
 FILLCELL_X1 FILLER_20_81 ();
 FILLCELL_X8 FILLER_20_85 ();
 FILLCELL_X1 FILLER_20_9 ();
 FILLCELL_X8 FILLER_20_95 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X1 FILLER_21_103 ();
 FILLCELL_X1 FILLER_21_104 ();
 FILLCELL_X1 FILLER_21_108 ();
 FILLCELL_X1 FILLER_21_109 ();
 FILLCELL_X8 FILLER_21_113 ();
 FILLCELL_X1 FILLER_21_121 ();
 FILLCELL_X8 FILLER_21_124 ();
 FILLCELL_X1 FILLER_21_132 ();
 FILLCELL_X1 FILLER_21_133 ();
 FILLCELL_X1 FILLER_21_136 ();
 FILLCELL_X1 FILLER_21_137 ();
 FILLCELL_X1 FILLER_21_138 ();
 FILLCELL_X1 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_15 ();
 FILLCELL_X8 FILLER_21_155 ();
 FILLCELL_X4 FILLER_21_163 ();
 FILLCELL_X1 FILLER_21_167 ();
 FILLCELL_X1 FILLER_21_171 ();
 FILLCELL_X1 FILLER_21_172 ();
 FILLCELL_X8 FILLER_21_189 ();
 FILLCELL_X1 FILLER_21_197 ();
 FILLCELL_X1 FILLER_21_198 ();
 FILLCELL_X1 FILLER_21_2 ();
 FILLCELL_X1 FILLER_21_20 ();
 FILLCELL_X32 FILLER_21_201 ();
 FILLCELL_X1 FILLER_21_21 ();
 FILLCELL_X1 FILLER_21_22 ();
 FILLCELL_X8 FILLER_21_233 ();
 FILLCELL_X4 FILLER_21_241 ();
 FILLCELL_X1 FILLER_21_39 ();
 FILLCELL_X1 FILLER_21_40 ();
 FILLCELL_X16 FILLER_21_43 ();
 FILLCELL_X4 FILLER_21_59 ();
 FILLCELL_X1 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_64 ();
 FILLCELL_X4 FILLER_21_68 ();
 FILLCELL_X1 FILLER_21_72 ();
 FILLCELL_X1 FILLER_21_73 ();
 FILLCELL_X1 FILLER_21_74 ();
 FILLCELL_X1 FILLER_21_77 ();
 FILLCELL_X1 FILLER_21_78 ();
 FILLCELL_X1 FILLER_21_8 ();
 FILLCELL_X1 FILLER_21_9 ();
 FILLCELL_X8 FILLER_21_95 ();
 FILLCELL_X1 FILLER_22_1 ();
 FILLCELL_X16 FILLER_22_121 ();
 FILLCELL_X8 FILLER_22_13 ();
 FILLCELL_X32 FILLER_22_147 ();
 FILLCELL_X32 FILLER_22_179 ();
 FILLCELL_X1 FILLER_22_2 ();
 FILLCELL_X4 FILLER_22_21 ();
 FILLCELL_X32 FILLER_22_211 ();
 FILLCELL_X1 FILLER_22_243 ();
 FILLCELL_X1 FILLER_22_244 ();
 FILLCELL_X1 FILLER_22_25 ();
 FILLCELL_X1 FILLER_22_29 ();
 FILLCELL_X1 FILLER_22_30 ();
 FILLCELL_X32 FILLER_22_34 ();
 FILLCELL_X16 FILLER_22_66 ();
 FILLCELL_X1 FILLER_22_7 ();
 FILLCELL_X1 FILLER_22_8 ();
 FILLCELL_X4 FILLER_22_82 ();
 FILLCELL_X32 FILLER_22_89 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_129 ();
 FILLCELL_X32 FILLER_23_161 ();
 FILLCELL_X32 FILLER_23_193 ();
 FILLCELL_X16 FILLER_23_225 ();
 FILLCELL_X4 FILLER_23_241 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X32 FILLER_23_97 ();
 FILLCELL_X8 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_105 ();
 FILLCELL_X1 FILLER_2_106 ();
 FILLCELL_X1 FILLER_2_110 ();
 FILLCELL_X1 FILLER_2_111 ();
 FILLCELL_X32 FILLER_2_115 ();
 FILLCELL_X1 FILLER_2_13 ();
 FILLCELL_X1 FILLER_2_14 ();
 FILLCELL_X1 FILLER_2_147 ();
 FILLCELL_X1 FILLER_2_15 ();
 FILLCELL_X4 FILLER_2_153 ();
 FILLCELL_X1 FILLER_2_157 ();
 FILLCELL_X1 FILLER_2_158 ();
 FILLCELL_X1 FILLER_2_159 ();
 FILLCELL_X4 FILLER_2_163 ();
 FILLCELL_X16 FILLER_2_170 ();
 FILLCELL_X4 FILLER_2_186 ();
 FILLCELL_X1 FILLER_2_19 ();
 FILLCELL_X1 FILLER_2_190 ();
 FILLCELL_X1 FILLER_2_191 ();
 FILLCELL_X1 FILLER_2_192 ();
 FILLCELL_X1 FILLER_2_197 ();
 FILLCELL_X1 FILLER_2_198 ();
 FILLCELL_X1 FILLER_2_20 ();
 FILLCELL_X16 FILLER_2_202 ();
 FILLCELL_X1 FILLER_2_221 ();
 FILLCELL_X1 FILLER_2_222 ();
 FILLCELL_X1 FILLER_2_226 ();
 FILLCELL_X1 FILLER_2_227 ();
 FILLCELL_X4 FILLER_2_231 ();
 FILLCELL_X1 FILLER_2_238 ();
 FILLCELL_X1 FILLER_2_239 ();
 FILLCELL_X1 FILLER_2_24 ();
 FILLCELL_X1 FILLER_2_243 ();
 FILLCELL_X1 FILLER_2_244 ();
 FILLCELL_X1 FILLER_2_25 ();
 FILLCELL_X1 FILLER_2_31 ();
 FILLCELL_X1 FILLER_2_32 ();
 FILLCELL_X8 FILLER_2_38 ();
 FILLCELL_X4 FILLER_2_46 ();
 FILLCELL_X1 FILLER_2_50 ();
 FILLCELL_X1 FILLER_2_51 ();
 FILLCELL_X1 FILLER_2_57 ();
 FILLCELL_X1 FILLER_2_58 ();
 FILLCELL_X16 FILLER_2_64 ();
 FILLCELL_X8 FILLER_2_80 ();
 FILLCELL_X4 FILLER_2_88 ();
 FILLCELL_X4 FILLER_2_9 ();
 FILLCELL_X1 FILLER_2_92 ();
 FILLCELL_X1 FILLER_2_98 ();
 FILLCELL_X1 FILLER_2_99 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_100 ();
 FILLCELL_X1 FILLER_3_104 ();
 FILLCELL_X1 FILLER_3_105 ();
 FILLCELL_X4 FILLER_3_108 ();
 FILLCELL_X1 FILLER_3_112 ();
 FILLCELL_X1 FILLER_3_116 ();
 FILLCELL_X1 FILLER_3_117 ();
 FILLCELL_X1 FILLER_3_121 ();
 FILLCELL_X1 FILLER_3_122 ();
 FILLCELL_X16 FILLER_3_126 ();
 FILLCELL_X8 FILLER_3_142 ();
 FILLCELL_X1 FILLER_3_150 ();
 FILLCELL_X1 FILLER_3_154 ();
 FILLCELL_X1 FILLER_3_155 ();
 FILLCELL_X1 FILLER_3_160 ();
 FILLCELL_X1 FILLER_3_161 ();
 FILLCELL_X1 FILLER_3_166 ();
 FILLCELL_X1 FILLER_3_167 ();
 FILLCELL_X8 FILLER_3_17 ();
 FILLCELL_X16 FILLER_3_170 ();
 FILLCELL_X4 FILLER_3_186 ();
 FILLCELL_X1 FILLER_3_190 ();
 FILLCELL_X1 FILLER_3_191 ();
 FILLCELL_X1 FILLER_3_192 ();
 FILLCELL_X1 FILLER_3_195 ();
 FILLCELL_X1 FILLER_3_196 ();
 FILLCELL_X1 FILLER_3_200 ();
 FILLCELL_X1 FILLER_3_201 ();
 FILLCELL_X1 FILLER_3_205 ();
 FILLCELL_X1 FILLER_3_206 ();
 FILLCELL_X8 FILLER_3_210 ();
 FILLCELL_X1 FILLER_3_220 ();
 FILLCELL_X1 FILLER_3_221 ();
 FILLCELL_X1 FILLER_3_222 ();
 FILLCELL_X8 FILLER_3_225 ();
 FILLCELL_X4 FILLER_3_233 ();
 FILLCELL_X1 FILLER_3_237 ();
 FILLCELL_X1 FILLER_3_238 ();
 FILLCELL_X1 FILLER_3_239 ();
 FILLCELL_X1 FILLER_3_243 ();
 FILLCELL_X1 FILLER_3_244 ();
 FILLCELL_X4 FILLER_3_25 ();
 FILLCELL_X1 FILLER_3_34 ();
 FILLCELL_X1 FILLER_3_35 ();
 FILLCELL_X8 FILLER_3_39 ();
 FILLCELL_X1 FILLER_3_47 ();
 FILLCELL_X1 FILLER_3_48 ();
 FILLCELL_X1 FILLER_3_49 ();
 FILLCELL_X1 FILLER_3_53 ();
 FILLCELL_X1 FILLER_3_54 ();
 FILLCELL_X1 FILLER_3_55 ();
 FILLCELL_X32 FILLER_3_59 ();
 FILLCELL_X8 FILLER_3_91 ();
 FILLCELL_X1 FILLER_3_99 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X1 FILLER_4_101 ();
 FILLCELL_X1 FILLER_4_106 ();
 FILLCELL_X1 FILLER_4_107 ();
 FILLCELL_X32 FILLER_4_111 ();
 FILLCELL_X32 FILLER_4_143 ();
 FILLCELL_X8 FILLER_4_175 ();
 FILLCELL_X1 FILLER_4_183 ();
 FILLCELL_X1 FILLER_4_184 ();
 FILLCELL_X1 FILLER_4_187 ();
 FILLCELL_X1 FILLER_4_188 ();
 FILLCELL_X1 FILLER_4_192 ();
 FILLCELL_X1 FILLER_4_193 ();
 FILLCELL_X1 FILLER_4_197 ();
 FILLCELL_X1 FILLER_4_198 ();
 FILLCELL_X32 FILLER_4_202 ();
 FILLCELL_X8 FILLER_4_234 ();
 FILLCELL_X1 FILLER_4_242 ();
 FILLCELL_X1 FILLER_4_243 ();
 FILLCELL_X1 FILLER_4_244 ();
 FILLCELL_X4 FILLER_4_33 ();
 FILLCELL_X1 FILLER_4_37 ();
 FILLCELL_X1 FILLER_4_38 ();
 FILLCELL_X1 FILLER_4_44 ();
 FILLCELL_X1 FILLER_4_45 ();
 FILLCELL_X1 FILLER_4_51 ();
 FILLCELL_X1 FILLER_4_52 ();
 FILLCELL_X1 FILLER_4_53 ();
 FILLCELL_X32 FILLER_4_57 ();
 FILLCELL_X8 FILLER_4_89 ();
 FILLCELL_X4 FILLER_4_97 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X4 FILLER_5_105 ();
 FILLCELL_X4 FILLER_5_112 ();
 FILLCELL_X1 FILLER_5_116 ();
 FILLCELL_X1 FILLER_5_117 ();
 FILLCELL_X1 FILLER_5_118 ();
 FILLCELL_X32 FILLER_5_123 ();
 FILLCELL_X16 FILLER_5_155 ();
 FILLCELL_X1 FILLER_5_171 ();
 FILLCELL_X1 FILLER_5_172 ();
 FILLCELL_X1 FILLER_5_173 ();
 FILLCELL_X32 FILLER_5_184 ();
 FILLCELL_X16 FILLER_5_216 ();
 FILLCELL_X8 FILLER_5_232 ();
 FILLCELL_X4 FILLER_5_240 ();
 FILLCELL_X1 FILLER_5_244 ();
 FILLCELL_X8 FILLER_5_33 ();
 FILLCELL_X4 FILLER_5_45 ();
 FILLCELL_X1 FILLER_5_49 ();
 FILLCELL_X1 FILLER_5_50 ();
 FILLCELL_X1 FILLER_5_51 ();
 FILLCELL_X32 FILLER_5_55 ();
 FILLCELL_X8 FILLER_5_87 ();
 FILLCELL_X8 FILLER_5_97 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X4 FILLER_6_100 ();
 FILLCELL_X1 FILLER_6_104 ();
 FILLCELL_X1 FILLER_6_105 ();
 FILLCELL_X4 FILLER_6_109 ();
 FILLCELL_X1 FILLER_6_113 ();
 FILLCELL_X32 FILLER_6_117 ();
 FILLCELL_X32 FILLER_6_149 ();
 FILLCELL_X16 FILLER_6_181 ();
 FILLCELL_X8 FILLER_6_197 ();
 FILLCELL_X1 FILLER_6_205 ();
 FILLCELL_X1 FILLER_6_206 ();
 FILLCELL_X1 FILLER_6_207 ();
 FILLCELL_X1 FILLER_6_210 ();
 FILLCELL_X1 FILLER_6_211 ();
 FILLCELL_X1 FILLER_6_212 ();
 FILLCELL_X1 FILLER_6_216 ();
 FILLCELL_X1 FILLER_6_217 ();
 FILLCELL_X16 FILLER_6_221 ();
 FILLCELL_X1 FILLER_6_237 ();
 FILLCELL_X1 FILLER_6_238 ();
 FILLCELL_X1 FILLER_6_239 ();
 FILLCELL_X1 FILLER_6_243 ();
 FILLCELL_X1 FILLER_6_244 ();
 FILLCELL_X8 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_44 ();
 FILLCELL_X8 FILLER_6_76 ();
 FILLCELL_X4 FILLER_6_84 ();
 FILLCELL_X1 FILLER_6_88 ();
 FILLCELL_X8 FILLER_6_92 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X8 FILLER_7_110 ();
 FILLCELL_X4 FILLER_7_118 ();
 FILLCELL_X1 FILLER_7_122 ();
 FILLCELL_X1 FILLER_7_123 ();
 FILLCELL_X1 FILLER_7_124 ();
 FILLCELL_X1 FILLER_7_129 ();
 FILLCELL_X1 FILLER_7_130 ();
 FILLCELL_X16 FILLER_7_134 ();
 FILLCELL_X1 FILLER_7_150 ();
 FILLCELL_X1 FILLER_7_151 ();
 FILLCELL_X1 FILLER_7_152 ();
 FILLCELL_X32 FILLER_7_156 ();
 FILLCELL_X8 FILLER_7_188 ();
 FILLCELL_X4 FILLER_7_196 ();
 FILLCELL_X1 FILLER_7_200 ();
 FILLCELL_X1 FILLER_7_201 ();
 FILLCELL_X1 FILLER_7_202 ();
 FILLCELL_X1 FILLER_7_206 ();
 FILLCELL_X1 FILLER_7_207 ();
 FILLCELL_X1 FILLER_7_211 ();
 FILLCELL_X1 FILLER_7_212 ();
 FILLCELL_X4 FILLER_7_216 ();
 FILLCELL_X1 FILLER_7_220 ();
 FILLCELL_X1 FILLER_7_221 ();
 FILLCELL_X16 FILLER_7_226 ();
 FILLCELL_X1 FILLER_7_242 ();
 FILLCELL_X1 FILLER_7_243 ();
 FILLCELL_X1 FILLER_7_244 ();
 FILLCELL_X1 FILLER_7_33 ();
 FILLCELL_X1 FILLER_7_37 ();
 FILLCELL_X1 FILLER_7_38 ();
 FILLCELL_X1 FILLER_7_42 ();
 FILLCELL_X1 FILLER_7_43 ();
 FILLCELL_X32 FILLER_7_46 ();
 FILLCELL_X32 FILLER_7_78 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X1 FILLER_8_104 ();
 FILLCELL_X1 FILLER_8_105 ();
 FILLCELL_X1 FILLER_8_106 ();
 FILLCELL_X1 FILLER_8_110 ();
 FILLCELL_X1 FILLER_8_111 ();
 FILLCELL_X16 FILLER_8_115 ();
 FILLCELL_X8 FILLER_8_131 ();
 FILLCELL_X4 FILLER_8_139 ();
 FILLCELL_X1 FILLER_8_143 ();
 FILLCELL_X1 FILLER_8_144 ();
 FILLCELL_X1 FILLER_8_145 ();
 FILLCELL_X4 FILLER_8_149 ();
 FILLCELL_X1 FILLER_8_157 ();
 FILLCELL_X1 FILLER_8_158 ();
 FILLCELL_X1 FILLER_8_162 ();
 FILLCELL_X1 FILLER_8_163 ();
 FILLCELL_X32 FILLER_8_167 ();
 FILLCELL_X8 FILLER_8_17 ();
 FILLCELL_X4 FILLER_8_199 ();
 FILLCELL_X1 FILLER_8_203 ();
 FILLCELL_X1 FILLER_8_204 ();
 FILLCELL_X1 FILLER_8_205 ();
 FILLCELL_X1 FILLER_8_209 ();
 FILLCELL_X1 FILLER_8_210 ();
 FILLCELL_X1 FILLER_8_214 ();
 FILLCELL_X1 FILLER_8_215 ();
 FILLCELL_X16 FILLER_8_218 ();
 FILLCELL_X4 FILLER_8_234 ();
 FILLCELL_X1 FILLER_8_238 ();
 FILLCELL_X1 FILLER_8_239 ();
 FILLCELL_X1 FILLER_8_243 ();
 FILLCELL_X1 FILLER_8_244 ();
 FILLCELL_X4 FILLER_8_25 ();
 FILLCELL_X32 FILLER_8_32 ();
 FILLCELL_X8 FILLER_8_64 ();
 FILLCELL_X4 FILLER_8_72 ();
 FILLCELL_X1 FILLER_8_76 ();
 FILLCELL_X1 FILLER_8_77 ();
 FILLCELL_X1 FILLER_8_78 ();
 FILLCELL_X4 FILLER_8_82 ();
 FILLCELL_X1 FILLER_8_86 ();
 FILLCELL_X1 FILLER_8_91 ();
 FILLCELL_X1 FILLER_8_92 ();
 FILLCELL_X8 FILLER_8_96 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X4 FILLER_9_118 ();
 FILLCELL_X1 FILLER_9_122 ();
 FILLCELL_X16 FILLER_9_126 ();
 FILLCELL_X8 FILLER_9_142 ();
 FILLCELL_X1 FILLER_9_150 ();
 FILLCELL_X1 FILLER_9_151 ();
 FILLCELL_X1 FILLER_9_152 ();
 FILLCELL_X1 FILLER_9_157 ();
 FILLCELL_X1 FILLER_9_158 ();
 FILLCELL_X32 FILLER_9_161 ();
 FILLCELL_X4 FILLER_9_17 ();
 FILLCELL_X4 FILLER_9_193 ();
 FILLCELL_X32 FILLER_9_207 ();
 FILLCELL_X1 FILLER_9_21 ();
 FILLCELL_X4 FILLER_9_239 ();
 FILLCELL_X1 FILLER_9_243 ();
 FILLCELL_X1 FILLER_9_244 ();
 FILLCELL_X1 FILLER_9_32 ();
 FILLCELL_X1 FILLER_9_33 ();
 FILLCELL_X1 FILLER_9_37 ();
 FILLCELL_X1 FILLER_9_38 ();
 FILLCELL_X1 FILLER_9_39 ();
 FILLCELL_X1 FILLER_9_43 ();
 FILLCELL_X1 FILLER_9_44 ();
 FILLCELL_X4 FILLER_9_48 ();
 FILLCELL_X16 FILLER_9_54 ();
 FILLCELL_X8 FILLER_9_70 ();
 FILLCELL_X4 FILLER_9_78 ();
 FILLCELL_X1 FILLER_9_82 ();
 FILLCELL_X32 FILLER_9_86 ();
 TAPCELL_X1 PHY_0 ();
 TAPCELL_X1 PHY_1 ();
 TAPCELL_X1 PHY_10 ();
 TAPCELL_X1 PHY_11 ();
 TAPCELL_X1 PHY_12 ();
 TAPCELL_X1 PHY_13 ();
 TAPCELL_X1 PHY_14 ();
 TAPCELL_X1 PHY_15 ();
 TAPCELL_X1 PHY_16 ();
 TAPCELL_X1 PHY_17 ();
 TAPCELL_X1 PHY_18 ();
 TAPCELL_X1 PHY_19 ();
 TAPCELL_X1 PHY_2 ();
 TAPCELL_X1 PHY_20 ();
 TAPCELL_X1 PHY_21 ();
 TAPCELL_X1 PHY_22 ();
 TAPCELL_X1 PHY_23 ();
 TAPCELL_X1 PHY_24 ();
 TAPCELL_X1 PHY_25 ();
 TAPCELL_X1 PHY_26 ();
 TAPCELL_X1 PHY_27 ();
 TAPCELL_X1 PHY_28 ();
 TAPCELL_X1 PHY_29 ();
 TAPCELL_X1 PHY_3 ();
 TAPCELL_X1 PHY_30 ();
 TAPCELL_X1 PHY_31 ();
 TAPCELL_X1 PHY_32 ();
 TAPCELL_X1 PHY_33 ();
 TAPCELL_X1 PHY_34 ();
 TAPCELL_X1 PHY_35 ();
 TAPCELL_X1 PHY_36 ();
 TAPCELL_X1 PHY_37 ();
 TAPCELL_X1 PHY_38 ();
 TAPCELL_X1 PHY_39 ();
 TAPCELL_X1 PHY_4 ();
 TAPCELL_X1 PHY_40 ();
 TAPCELL_X1 PHY_41 ();
 TAPCELL_X1 PHY_42 ();
 TAPCELL_X1 PHY_43 ();
 TAPCELL_X1 PHY_44 ();
 TAPCELL_X1 PHY_45 ();
 TAPCELL_X1 PHY_46 ();
 TAPCELL_X1 PHY_47 ();
 TAPCELL_X1 PHY_5 ();
 TAPCELL_X1 PHY_6 ();
 TAPCELL_X1 PHY_7 ();
 TAPCELL_X1 PHY_8 ();
 TAPCELL_X1 PHY_9 ();
 INV_X4 _225_ (.A(net10),
    .ZN(_130_));
 NAND2_X1 _227_ (.A1(_130_),
    .A2(net9),
    .ZN(_132_));
 INV_X2 _228_ (.A(net12),
    .ZN(_000_));
 NAND2_X2 _229_ (.A1(_000_),
    .A2(net11),
    .ZN(_001_));
 NOR2_X1 _230_ (.A1(_132_),
    .A2(_001_),
    .ZN(_002_));
 INV_X1 _231_ (.A(_163_),
    .ZN(_003_));
 NAND2_X1 _232_ (.A1(_002_),
    .A2(_003_),
    .ZN(_004_));
 INV_X4 _233_ (.A(net9),
    .ZN(_005_));
 NAND2_X1 _234_ (.A1(_005_),
    .A2(net10),
    .ZN(_006_));
 NOR2_X2 _235_ (.A1(_006_),
    .A2(_001_),
    .ZN(_007_));
 NAND2_X1 _236_ (.A1(_007_),
    .A2(_206_),
    .ZN(_008_));
 NAND2_X1 _237_ (.A1(_004_),
    .A2(_008_),
    .ZN(_009_));
 NAND2_X1 _238_ (.A1(_130_),
    .A2(_005_),
    .ZN(_010_));
 NOR2_X2 _239_ (.A1(_010_),
    .A2(_001_),
    .ZN(_011_));
 INV_X1 _240_ (.A(net3),
    .ZN(_142_));
 NAND2_X1 _241_ (.A1(_011_),
    .A2(_142_),
    .ZN(_012_));
 INV_X2 _242_ (.A(net11),
    .ZN(_013_));
 NAND2_X1 _243_ (.A1(_013_),
    .A2(_000_),
    .ZN(_014_));
 NAND2_X1 _244_ (.A1(net10),
    .A2(net9),
    .ZN(_015_));
 NOR2_X1 _245_ (.A1(_014_),
    .A2(_015_),
    .ZN(_016_));
 INV_X1 _246_ (.A(_206_),
    .ZN(_017_));
 NAND2_X1 _247_ (.A1(_016_),
    .A2(_017_),
    .ZN(_018_));
 NAND2_X1 _248_ (.A1(_012_),
    .A2(_018_),
    .ZN(_019_));
 NOR2_X1 _249_ (.A1(_009_),
    .A2(_019_),
    .ZN(_020_));
 NOR2_X1 _250_ (.A1(_130_),
    .A2(net9),
    .ZN(_021_));
 NOR2_X2 _251_ (.A1(net11),
    .A2(net12),
    .ZN(_022_));
 NAND2_X1 _252_ (.A1(_021_),
    .A2(_022_),
    .ZN(_023_));
 INV_X1 _253_ (.A(_023_),
    .ZN(_024_));
 NAND2_X1 _254_ (.A1(_024_),
    .A2(_163_),
    .ZN(_025_));
 NOR2_X1 _255_ (.A1(_014_),
    .A2(_132_),
    .ZN(_026_));
 NAND2_X1 _256_ (.A1(_026_),
    .A2(_141_),
    .ZN(_027_));
 NAND2_X1 _257_ (.A1(_025_),
    .A2(_027_),
    .ZN(_028_));
 NOR2_X2 _258_ (.A1(net10),
    .A2(net9),
    .ZN(_029_));
 NAND2_X1 _259_ (.A1(_029_),
    .A2(_022_),
    .ZN(_030_));
 NOR2_X1 _260_ (.A1(_030_),
    .A2(_145_),
    .ZN(_031_));
 NOR2_X1 _261_ (.A1(_028_),
    .A2(_031_),
    .ZN(_032_));
 NAND2_X1 _262_ (.A1(_013_),
    .A2(net12),
    .ZN(_033_));
 INV_X2 _263_ (.A(_033_),
    .ZN(_034_));
 INV_X1 _264_ (.A(_195_),
    .ZN(_035_));
 NAND3_X1 _265_ (.A1(_034_),
    .A2(_029_),
    .A3(_035_),
    .ZN(_036_));
 NOR2_X2 _266_ (.A1(_013_),
    .A2(net12),
    .ZN(_037_));
 INV_X1 _267_ (.A(_015_),
    .ZN(_038_));
 NAND3_X1 _268_ (.A1(_037_),
    .A2(_038_),
    .A3(_195_),
    .ZN(_039_));
 NAND2_X1 _269_ (.A1(_036_),
    .A2(_039_),
    .ZN(_040_));
 NOR2_X2 _270_ (.A1(_005_),
    .A2(net10),
    .ZN(_041_));
 NAND2_X2 _271_ (.A1(_034_),
    .A2(_041_),
    .ZN(_042_));
 INV_X1 _272_ (.A(_194_),
    .ZN(_043_));
 NOR2_X1 _273_ (.A1(_042_),
    .A2(_043_),
    .ZN(_044_));
 NOR2_X1 _274_ (.A1(_040_),
    .A2(_044_),
    .ZN(_045_));
 NAND3_X1 _275_ (.A1(_020_),
    .A2(_032_),
    .A3(_045_),
    .ZN(net15));
 NAND2_X1 _276_ (.A1(net1),
    .A2(net8),
    .ZN(_046_));
 INV_X1 _277_ (.A(_046_),
    .ZN(_197_));
 NAND2_X1 _278_ (.A1(net7),
    .A2(net2),
    .ZN(_151_));
 NAND2_X1 _279_ (.A1(net5),
    .A2(net4),
    .ZN(_147_));
 NAND2_X1 _280_ (.A1(net3),
    .A2(net6),
    .ZN(_146_));
 NAND2_X1 _281_ (.A1(_007_),
    .A2(_202_),
    .ZN(_047_));
 INV_X1 _282_ (.A(_180_),
    .ZN(_048_));
 NAND2_X1 _283_ (.A1(_002_),
    .A2(_048_),
    .ZN(_049_));
 NAND2_X1 _284_ (.A1(_047_),
    .A2(_049_),
    .ZN(_050_));
 INV_X2 _285_ (.A(net4),
    .ZN(_154_));
 NAND2_X1 _286_ (.A1(_011_),
    .A2(_154_),
    .ZN(_051_));
 INV_X1 _287_ (.A(_202_),
    .ZN(_052_));
 NAND2_X1 _288_ (.A1(_016_),
    .A2(_052_),
    .ZN(_053_));
 NAND2_X1 _289_ (.A1(_051_),
    .A2(_053_),
    .ZN(_054_));
 NOR2_X1 _290_ (.A1(_050_),
    .A2(_054_),
    .ZN(_055_));
 NAND2_X1 _291_ (.A1(_024_),
    .A2(_180_),
    .ZN(_056_));
 NAND2_X1 _292_ (.A1(_026_),
    .A2(_157_),
    .ZN(_057_));
 NAND2_X1 _293_ (.A1(_056_),
    .A2(_057_),
    .ZN(_058_));
 NOR2_X1 _294_ (.A1(_030_),
    .A2(_160_),
    .ZN(_059_));
 NOR2_X1 _295_ (.A1(_058_),
    .A2(_059_),
    .ZN(_060_));
 INV_X1 _296_ (.A(_199_),
    .ZN(_061_));
 NAND3_X1 _297_ (.A1(_034_),
    .A2(_029_),
    .A3(_061_),
    .ZN(_062_));
 NAND3_X1 _298_ (.A1(_037_),
    .A2(_038_),
    .A3(_199_),
    .ZN(_063_));
 NAND2_X1 _299_ (.A1(_062_),
    .A2(_063_),
    .ZN(_064_));
 INV_X1 _300_ (.A(_198_),
    .ZN(_065_));
 NOR2_X1 _301_ (.A1(_042_),
    .A2(_065_),
    .ZN(_066_));
 NOR2_X1 _302_ (.A1(_064_),
    .A2(_066_),
    .ZN(_067_));
 NAND3_X1 _303_ (.A1(_055_),
    .A2(_060_),
    .A3(_067_),
    .ZN(net16));
 NAND2_X1 _304_ (.A1(net8),
    .A2(net2),
    .ZN(_068_));
 INV_X1 _305_ (.A(_068_),
    .ZN(_166_));
 NAND2_X1 _306_ (.A1(net4),
    .A2(net6),
    .ZN(_069_));
 INV_X1 _307_ (.A(_069_),
    .ZN(_200_));
 OR2_X1 _308_ (.A1(_030_),
    .A2(_159_),
    .ZN(_070_));
 NAND2_X1 _309_ (.A1(_026_),
    .A2(_156_),
    .ZN(_071_));
 NAND3_X1 _310_ (.A1(_034_),
    .A2(_041_),
    .A3(_169_),
    .ZN(_072_));
 NAND3_X1 _311_ (.A1(_070_),
    .A2(_071_),
    .A3(_072_),
    .ZN(net17));
 NAND2_X1 _312_ (.A1(net3),
    .A2(net8),
    .ZN(_175_));
 NAND2_X1 _313_ (.A1(net7),
    .A2(net4),
    .ZN(_073_));
 INV_X1 _314_ (.A(_073_),
    .ZN(_170_));
 NOR2_X1 _315_ (.A1(_042_),
    .A2(_178_),
    .ZN(net18));
 INV_X1 _316_ (.A(_182_),
    .ZN(_074_));
 NOR2_X1 _317_ (.A1(_042_),
    .A2(_074_),
    .ZN(net19));
 INV_X1 _318_ (.A(_181_),
    .ZN(_075_));
 NOR2_X1 _319_ (.A1(_042_),
    .A2(_075_),
    .ZN(net20));
 NOR2_X1 _320_ (.A1(_033_),
    .A2(_006_),
    .ZN(_076_));
 NOR2_X1 _321_ (.A1(_195_),
    .A2(_199_),
    .ZN(_077_));
 NOR2_X1 _322_ (.A1(_213_),
    .A2(_222_),
    .ZN(_078_));
 NAND2_X1 _323_ (.A1(_077_),
    .A2(_078_),
    .ZN(_079_));
 NAND2_X1 _324_ (.A1(_076_),
    .A2(_079_),
    .ZN(_080_));
 AOI21_X1 _325_ (.A(_203_),
    .B1(_061_),
    .B2(_207_),
    .ZN(_081_));
 NAND2_X1 _326_ (.A1(_077_),
    .A2(_139_),
    .ZN(_082_));
 NAND2_X1 _327_ (.A1(_081_),
    .A2(_082_),
    .ZN(_083_));
 NOR2_X1 _328_ (.A1(_080_),
    .A2(_083_),
    .ZN(_084_));
 INV_X1 _329_ (.A(_186_),
    .ZN(_085_));
 AOI21_X1 _330_ (.A(_085_),
    .B1(_042_),
    .B2(_023_),
    .ZN(_086_));
 NOR2_X1 _331_ (.A1(_084_),
    .A2(_086_),
    .ZN(_087_));
 NAND2_X1 _332_ (.A1(_002_),
    .A2(_085_),
    .ZN(_088_));
 INV_X1 _333_ (.A(_212_),
    .ZN(_089_));
 NAND2_X1 _334_ (.A1(_016_),
    .A2(_089_),
    .ZN(_090_));
 NAND2_X1 _335_ (.A1(_088_),
    .A2(_090_),
    .ZN(_091_));
 INV_X1 _336_ (.A(_213_),
    .ZN(_092_));
 NAND2_X1 _337_ (.A1(_037_),
    .A2(_038_),
    .ZN(_093_));
 NAND2_X1 _338_ (.A1(_022_),
    .A2(_130_),
    .ZN(_094_));
 AOI21_X1 _339_ (.A(_092_),
    .B1(_093_),
    .B2(_094_),
    .ZN(_095_));
 NOR2_X1 _340_ (.A1(_091_),
    .A2(_095_),
    .ZN(_096_));
 INV_X1 _341_ (.A(net1),
    .ZN(_210_));
 NAND2_X1 _342_ (.A1(_011_),
    .A2(_210_),
    .ZN(_097_));
 NAND2_X1 _343_ (.A1(_007_),
    .A2(_212_),
    .ZN(_098_));
 NAND2_X1 _344_ (.A1(_097_),
    .A2(_098_),
    .ZN(_099_));
 NOR3_X1 _345_ (.A1(_010_),
    .A2(_033_),
    .A3(_213_),
    .ZN(_100_));
 NOR2_X1 _346_ (.A1(_099_),
    .A2(_100_),
    .ZN(_101_));
 NAND3_X1 _347_ (.A1(_087_),
    .A2(_096_),
    .A3(_101_),
    .ZN(net13));
 NAND2_X1 _348_ (.A1(net5),
    .A2(net2),
    .ZN(_102_));
 INV_X1 _349_ (.A(_102_),
    .ZN(_217_));
 INV_X1 _350_ (.A(_189_),
    .ZN(_135_));
 INV_X1 _351_ (.A(_083_),
    .ZN(_103_));
 NOR2_X1 _352_ (.A1(_103_),
    .A2(_080_),
    .ZN(_104_));
 NAND2_X1 _353_ (.A1(_041_),
    .A2(_037_),
    .ZN(_105_));
 NAND2_X1 _354_ (.A1(_105_),
    .A2(_135_),
    .ZN(_106_));
 NAND2_X1 _355_ (.A1(_023_),
    .A2(_189_),
    .ZN(_107_));
 NAND2_X1 _356_ (.A1(_106_),
    .A2(_107_),
    .ZN(_108_));
 INV_X1 _357_ (.A(_108_),
    .ZN(_109_));
 NOR2_X1 _358_ (.A1(_104_),
    .A2(_109_),
    .ZN(_110_));
 INV_X1 _359_ (.A(_221_),
    .ZN(_111_));
 NAND2_X1 _360_ (.A1(_016_),
    .A2(_111_),
    .ZN(_112_));
 NAND3_X1 _361_ (.A1(_037_),
    .A2(_038_),
    .A3(_222_),
    .ZN(_113_));
 NAND2_X1 _362_ (.A1(_112_),
    .A2(_113_),
    .ZN(_114_));
 NAND3_X1 _363_ (.A1(_034_),
    .A2(_041_),
    .A3(_219_),
    .ZN(_115_));
 INV_X1 _364_ (.A(_222_),
    .ZN(_116_));
 NAND3_X1 _365_ (.A1(_034_),
    .A2(_029_),
    .A3(_116_),
    .ZN(_117_));
 NAND2_X1 _366_ (.A1(_115_),
    .A2(_117_),
    .ZN(_118_));
 NOR2_X1 _367_ (.A1(_114_),
    .A2(_118_),
    .ZN(_119_));
 INV_X1 _368_ (.A(net2),
    .ZN(_220_));
 NAND2_X1 _369_ (.A1(_011_),
    .A2(_220_),
    .ZN(_120_));
 NAND2_X1 _370_ (.A1(_007_),
    .A2(_221_),
    .ZN(_121_));
 NAND2_X1 _371_ (.A1(_120_),
    .A2(_121_),
    .ZN(_122_));
 NAND3_X1 _372_ (.A1(_029_),
    .A2(_022_),
    .A3(_188_),
    .ZN(_123_));
 NAND3_X1 _373_ (.A1(_041_),
    .A2(_022_),
    .A3(_185_),
    .ZN(_124_));
 NAND2_X1 _374_ (.A1(_123_),
    .A2(_124_),
    .ZN(_125_));
 NOR2_X1 _375_ (.A1(_122_),
    .A2(_125_),
    .ZN(_126_));
 NAND3_X1 _376_ (.A1(_110_),
    .A2(_119_),
    .A3(_126_),
    .ZN(net14));
 NAND2_X1 _377_ (.A1(net5),
    .A2(net3),
    .ZN(_133_));
 INV_X1 _378_ (.A(_173_),
    .ZN(_176_));
 INV_X1 _379_ (.A(_140_),
    .ZN(_155_));
 INV_X1 _380_ (.A(_168_),
    .ZN(_174_));
 INV_X1 _381_ (.A(_187_),
    .ZN(_143_));
 NAND2_X1 _382_ (.A1(net7),
    .A2(net1),
    .ZN(_127_));
 INV_X1 _383_ (.A(_127_),
    .ZN(_191_));
 INV_X1 _384_ (.A(_153_),
    .ZN(_196_));
 INV_X1 _385_ (.A(_177_),
    .ZN(_179_));
 INV_X1 _386_ (.A(_214_),
    .ZN(_184_));
 INV_X1 _387_ (.A(_137_),
    .ZN(_192_));
 INV_X1 _388_ (.A(_148_),
    .ZN(_201_));
 INV_X1 _389_ (.A(_152_),
    .ZN(_162_));
 INV_X1 _390_ (.A(net8),
    .ZN(_158_));
 INV_X2 _391_ (.A(net7),
    .ZN(_138_));
 INV_X1 _392_ (.A(net5),
    .ZN(_211_));
 NAND2_X1 _393_ (.A1(net1),
    .A2(net6),
    .ZN(_128_));
 INV_X1 _394_ (.A(_128_),
    .ZN(_218_));
 INV_X1 _395_ (.A(net6),
    .ZN(_183_));
 INV_X1 _396_ (.A(_193_),
    .ZN(_150_));
 INV_X1 _397_ (.A(_190_),
    .ZN(_134_));
 FA_X1 _398_ (.A(_133_),
    .B(_134_),
    .CI(_135_),
    .CO(_136_),
    .S(_137_));
 FA_X1 _399_ (.A(net3),
    .B(_138_),
    .CI(_139_),
    .CO(_140_),
    .S(_141_));
 FA_X1 _400_ (.A(_142_),
    .B(_138_),
    .CI(_143_),
    .CO(_144_),
    .S(_145_));
 FA_X1 _401_ (.A(_136_),
    .B(_146_),
    .CI(_147_),
    .CO(_148_),
    .S(_149_));
 FA_X1 _402_ (.A(_150_),
    .B(_151_),
    .CI(_149_),
    .CO(_152_),
    .S(_153_));
 FA_X1 _403_ (.A(_154_),
    .B(net8),
    .CI(_155_),
    .CO(_156_),
    .S(_157_));
 FA_X1 _404_ (.A(_154_),
    .B(_158_),
    .CI(_144_),
    .CO(_159_),
    .S(_160_));
 FA_X1 _405_ (.A(_161_),
    .B(_162_),
    .CI(_163_),
    .CO(_164_),
    .S(_165_));
 FA_X1 _406_ (.A(_166_),
    .B(_165_),
    .CI(_167_),
    .CO(_168_),
    .S(_169_));
 FA_X1 _407_ (.A(_170_),
    .B(_171_),
    .CI(_164_),
    .CO(_172_),
    .S(_173_));
 FA_X1 _408_ (.A(_174_),
    .B(_175_),
    .CI(_176_),
    .CO(_177_),
    .S(_178_));
 FA_X1 _409_ (.A(_179_),
    .B(_180_),
    .CI(_172_),
    .CO(_181_),
    .S(_182_));
 FA_X1 _410_ (.A(net2),
    .B(_183_),
    .CI(_184_),
    .CO(_139_),
    .S(_185_));
 FA_X1 _411_ (.A(net2),
    .B(net6),
    .CI(_186_),
    .CO(_187_),
    .S(_188_));
 HA_X1 _412_ (.A(_191_),
    .B(_192_),
    .CO(_193_),
    .S(_194_));
 HA_X1 _413_ (.A(_196_),
    .B(_197_),
    .CO(_167_),
    .S(_198_));
 HA_X1 _414_ (.A(_200_),
    .B(_201_),
    .CO(_171_),
    .S(_161_));
 HA_X1 _415_ (.A(_154_),
    .B(_158_),
    .CO(_202_),
    .S(_199_));
 HA_X1 _416_ (.A(net4),
    .B(_158_),
    .CO(_203_),
    .S(_204_));
 HA_X1 _417_ (.A(net4),
    .B(net8),
    .CO(_180_),
    .S(_205_));
 HA_X1 _418_ (.A(_142_),
    .B(_138_),
    .CO(_206_),
    .S(_195_));
 HA_X1 _419_ (.A(net3),
    .B(_138_),
    .CO(_207_),
    .S(_208_));
 HA_X1 _420_ (.A(net3),
    .B(net7),
    .CO(_163_),
    .S(_209_));
 HA_X1 _421_ (.A(_210_),
    .B(_211_),
    .CO(_212_),
    .S(_213_));
 HA_X1 _422_ (.A(_210_),
    .B(net5),
    .CO(_214_),
    .S(_215_));
 HA_X1 _423_ (.A(net1),
    .B(net5),
    .CO(_186_),
    .S(_216_));
 HA_X1 _424_ (.A(_217_),
    .B(_218_),
    .CO(_190_),
    .S(_219_));
 HA_X1 _425_ (.A(_220_),
    .B(_183_),
    .CO(_221_),
    .S(_222_));
 HA_X1 _426_ (.A(net2),
    .B(net6),
    .CO(_189_),
    .S(_223_));
 CLKBUF_X2 input1 (.A(A[0]),
    .Z(net1));
 BUF_X2 input10 (.A(CTRL[1]),
    .Z(net10));
 BUF_X1 input11 (.A(CTRL[2]),
    .Z(net11));
 CLKBUF_X2 input12 (.A(CTRL[3]),
    .Z(net12));
 CLKBUF_X3 input2 (.A(A[1]),
    .Z(net2));
 CLKBUF_X3 input3 (.A(A[2]),
    .Z(net3));
 BUF_X2 input4 (.A(A[3]),
    .Z(net4));
 BUF_X2 input5 (.A(B[0]),
    .Z(net5));
 BUF_X2 input6 (.A(B[1]),
    .Z(net6));
 BUF_X2 input7 (.A(B[2]),
    .Z(net7));
 BUF_X2 input8 (.A(B[3]),
    .Z(net8));
 BUF_X2 input9 (.A(CTRL[0]),
    .Z(net9));
 BUF_X1 output13 (.A(net13),
    .Z(Y[0]));
 BUF_X1 output14 (.A(net14),
    .Z(Y[1]));
 BUF_X1 output15 (.A(net15),
    .Z(Y[2]));
 BUF_X1 output16 (.A(net16),
    .Z(Y[3]));
 BUF_X1 output17 (.A(net17),
    .Z(Y[4]));
 BUF_X1 output18 (.A(net18),
    .Z(Y[5]));
 BUF_X1 output19 (.A(net19),
    .Z(Y[6]));
 BUF_X1 output20 (.A(net20),
    .Z(Y[7]));
endmodule

module alu_4 (A,
    B,
    CTRL,
    Y);
 input [3:0] A;
 input [3:0] B;
 input [3:0] CTRL;
 output [7:0] Y;

 wire VDD;
 wire VSS;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _107_;
 wire _109_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 FILLCELL_X16 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_100 ();
 FILLCELL_X32 FILLER_0_132 ();
 FILLCELL_X32 FILLER_0_164 ();
 FILLCELL_X1 FILLER_0_17 ();
 FILLCELL_X1 FILLER_0_18 ();
 FILLCELL_X32 FILLER_0_196 ();
 FILLCELL_X16 FILLER_0_228 ();
 FILLCELL_X1 FILLER_0_23 ();
 FILLCELL_X1 FILLER_0_24 ();
 FILLCELL_X1 FILLER_0_244 ();
 FILLCELL_X1 FILLER_0_30 ();
 FILLCELL_X1 FILLER_0_31 ();
 FILLCELL_X32 FILLER_0_36 ();
 FILLCELL_X32 FILLER_0_68 ();
 FILLCELL_X16 FILLER_10_1 ();
 FILLCELL_X8 FILLER_10_100 ();
 FILLCELL_X4 FILLER_10_108 ();
 FILLCELL_X1 FILLER_10_112 ();
 FILLCELL_X1 FILLER_10_113 ();
 FILLCELL_X1 FILLER_10_114 ();
 FILLCELL_X8 FILLER_10_119 ();
 FILLCELL_X1 FILLER_10_127 ();
 FILLCELL_X1 FILLER_10_128 ();
 FILLCELL_X32 FILLER_10_133 ();
 FILLCELL_X16 FILLER_10_165 ();
 FILLCELL_X4 FILLER_10_17 ();
 FILLCELL_X8 FILLER_10_181 ();
 FILLCELL_X4 FILLER_10_189 ();
 FILLCELL_X1 FILLER_10_193 ();
 FILLCELL_X1 FILLER_10_194 ();
 FILLCELL_X32 FILLER_10_197 ();
 FILLCELL_X1 FILLER_10_21 ();
 FILLCELL_X1 FILLER_10_22 ();
 FILLCELL_X16 FILLER_10_229 ();
 FILLCELL_X4 FILLER_10_27 ();
 FILLCELL_X1 FILLER_10_31 ();
 FILLCELL_X1 FILLER_10_32 ();
 FILLCELL_X1 FILLER_10_43 ();
 FILLCELL_X1 FILLER_10_44 ();
 FILLCELL_X1 FILLER_10_49 ();
 FILLCELL_X1 FILLER_10_50 ();
 FILLCELL_X16 FILLER_10_54 ();
 FILLCELL_X8 FILLER_10_70 ();
 FILLCELL_X4 FILLER_10_78 ();
 FILLCELL_X8 FILLER_10_84 ();
 FILLCELL_X4 FILLER_10_92 ();
 FILLCELL_X1 FILLER_10_96 ();
 FILLCELL_X1 FILLER_10_97 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_107 ();
 FILLCELL_X4 FILLER_11_139 ();
 FILLCELL_X1 FILLER_11_143 ();
 FILLCELL_X1 FILLER_11_144 ();
 FILLCELL_X32 FILLER_11_149 ();
 FILLCELL_X32 FILLER_11_181 ();
 FILLCELL_X1 FILLER_11_213 ();
 FILLCELL_X1 FILLER_11_214 ();
 FILLCELL_X1 FILLER_11_215 ();
 FILLCELL_X1 FILLER_11_220 ();
 FILLCELL_X1 FILLER_11_221 ();
 FILLCELL_X16 FILLER_11_225 ();
 FILLCELL_X4 FILLER_11_241 ();
 FILLCELL_X4 FILLER_11_33 ();
 FILLCELL_X1 FILLER_11_37 ();
 FILLCELL_X1 FILLER_11_38 ();
 FILLCELL_X32 FILLER_11_43 ();
 FILLCELL_X32 FILLER_11_75 ();
 FILLCELL_X16 FILLER_12_1 ();
 FILLCELL_X1 FILLER_12_102 ();
 FILLCELL_X1 FILLER_12_103 ();
 FILLCELL_X1 FILLER_12_104 ();
 FILLCELL_X32 FILLER_12_108 ();
 FILLCELL_X16 FILLER_12_140 ();
 FILLCELL_X1 FILLER_12_159 ();
 FILLCELL_X1 FILLER_12_160 ();
 FILLCELL_X32 FILLER_12_164 ();
 FILLCELL_X8 FILLER_12_17 ();
 FILLCELL_X8 FILLER_12_196 ();
 FILLCELL_X1 FILLER_12_204 ();
 FILLCELL_X1 FILLER_12_205 ();
 FILLCELL_X1 FILLER_12_206 ();
 FILLCELL_X4 FILLER_12_210 ();
 FILLCELL_X1 FILLER_12_217 ();
 FILLCELL_X1 FILLER_12_218 ();
 FILLCELL_X16 FILLER_12_222 ();
 FILLCELL_X1 FILLER_12_238 ();
 FILLCELL_X1 FILLER_12_239 ();
 FILLCELL_X1 FILLER_12_243 ();
 FILLCELL_X1 FILLER_12_244 ();
 FILLCELL_X4 FILLER_12_25 ();
 FILLCELL_X1 FILLER_12_29 ();
 FILLCELL_X1 FILLER_12_30 ();
 FILLCELL_X1 FILLER_12_31 ();
 FILLCELL_X32 FILLER_12_34 ();
 FILLCELL_X32 FILLER_12_66 ();
 FILLCELL_X4 FILLER_12_98 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X4 FILLER_13_102 ();
 FILLCELL_X1 FILLER_13_109 ();
 FILLCELL_X1 FILLER_13_110 ();
 FILLCELL_X16 FILLER_13_114 ();
 FILLCELL_X8 FILLER_13_130 ();
 FILLCELL_X4 FILLER_13_138 ();
 FILLCELL_X1 FILLER_13_158 ();
 FILLCELL_X1 FILLER_13_159 ();
 FILLCELL_X1 FILLER_13_163 ();
 FILLCELL_X1 FILLER_13_164 ();
 FILLCELL_X16 FILLER_13_167 ();
 FILLCELL_X8 FILLER_13_183 ();
 FILLCELL_X4 FILLER_13_191 ();
 FILLCELL_X1 FILLER_13_195 ();
 FILLCELL_X1 FILLER_13_196 ();
 FILLCELL_X1 FILLER_13_197 ();
 FILLCELL_X1 FILLER_13_214 ();
 FILLCELL_X1 FILLER_13_215 ();
 FILLCELL_X1 FILLER_13_219 ();
 FILLCELL_X1 FILLER_13_220 ();
 FILLCELL_X16 FILLER_13_223 ();
 FILLCELL_X4 FILLER_13_239 ();
 FILLCELL_X1 FILLER_13_243 ();
 FILLCELL_X1 FILLER_13_244 ();
 FILLCELL_X4 FILLER_13_33 ();
 FILLCELL_X1 FILLER_13_37 ();
 FILLCELL_X1 FILLER_13_38 ();
 FILLCELL_X32 FILLER_13_41 ();
 FILLCELL_X8 FILLER_13_73 ();
 FILLCELL_X1 FILLER_13_81 ();
 FILLCELL_X1 FILLER_13_82 ();
 FILLCELL_X1 FILLER_13_83 ();
 FILLCELL_X16 FILLER_13_86 ();
 FILLCELL_X16 FILLER_14_1 ();
 FILLCELL_X1 FILLER_14_116 ();
 FILLCELL_X1 FILLER_14_117 ();
 FILLCELL_X16 FILLER_14_120 ();
 FILLCELL_X1 FILLER_14_136 ();
 FILLCELL_X1 FILLER_14_137 ();
 FILLCELL_X1 FILLER_14_138 ();
 FILLCELL_X1 FILLER_14_155 ();
 FILLCELL_X1 FILLER_14_156 ();
 FILLCELL_X32 FILLER_14_159 ();
 FILLCELL_X4 FILLER_14_17 ();
 FILLCELL_X1 FILLER_14_193 ();
 FILLCELL_X1 FILLER_14_194 ();
 FILLCELL_X1 FILLER_14_211 ();
 FILLCELL_X1 FILLER_14_212 ();
 FILLCELL_X16 FILLER_14_215 ();
 FILLCELL_X4 FILLER_14_23 ();
 FILLCELL_X8 FILLER_14_231 ();
 FILLCELL_X4 FILLER_14_239 ();
 FILLCELL_X1 FILLER_14_243 ();
 FILLCELL_X1 FILLER_14_244 ();
 FILLCELL_X1 FILLER_14_37 ();
 FILLCELL_X1 FILLER_14_38 ();
 FILLCELL_X1 FILLER_14_39 ();
 FILLCELL_X16 FILLER_14_42 ();
 FILLCELL_X8 FILLER_14_58 ();
 FILLCELL_X4 FILLER_14_66 ();
 FILLCELL_X1 FILLER_14_80 ();
 FILLCELL_X1 FILLER_14_81 ();
 FILLCELL_X1 FILLER_14_98 ();
 FILLCELL_X1 FILLER_14_99 ();
 FILLCELL_X8 FILLER_15_1 ();
 FILLCELL_X1 FILLER_15_10 ();
 FILLCELL_X16 FILLER_15_120 ();
 FILLCELL_X1 FILLER_15_13 ();
 FILLCELL_X8 FILLER_15_136 ();
 FILLCELL_X1 FILLER_15_14 ();
 FILLCELL_X4 FILLER_15_144 ();
 FILLCELL_X1 FILLER_15_148 ();
 FILLCELL_X32 FILLER_15_151 ();
 FILLCELL_X1 FILLER_15_18 ();
 FILLCELL_X32 FILLER_15_183 ();
 FILLCELL_X1 FILLER_15_19 ();
 FILLCELL_X16 FILLER_15_215 ();
 FILLCELL_X8 FILLER_15_231 ();
 FILLCELL_X4 FILLER_15_239 ();
 FILLCELL_X1 FILLER_15_243 ();
 FILLCELL_X1 FILLER_15_244 ();
 FILLCELL_X32 FILLER_15_30 ();
 FILLCELL_X8 FILLER_15_62 ();
 FILLCELL_X4 FILLER_15_70 ();
 FILLCELL_X1 FILLER_15_76 ();
 FILLCELL_X1 FILLER_15_77 ();
 FILLCELL_X32 FILLER_15_88 ();
 FILLCELL_X1 FILLER_15_9 ();
 FILLCELL_X16 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_106 ();
 FILLCELL_X32 FILLER_16_138 ();
 FILLCELL_X1 FILLER_16_17 ();
 FILLCELL_X16 FILLER_16_170 ();
 FILLCELL_X1 FILLER_16_18 ();
 FILLCELL_X1 FILLER_16_186 ();
 FILLCELL_X1 FILLER_16_187 ();
 FILLCELL_X1 FILLER_16_19 ();
 FILLCELL_X32 FILLER_16_191 ();
 FILLCELL_X16 FILLER_16_223 ();
 FILLCELL_X8 FILLER_16_23 ();
 FILLCELL_X4 FILLER_16_239 ();
 FILLCELL_X1 FILLER_16_243 ();
 FILLCELL_X1 FILLER_16_244 ();
 FILLCELL_X4 FILLER_16_31 ();
 FILLCELL_X1 FILLER_16_38 ();
 FILLCELL_X1 FILLER_16_39 ();
 FILLCELL_X32 FILLER_16_42 ();
 FILLCELL_X32 FILLER_16_74 ();
 FILLCELL_X16 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_110 ();
 FILLCELL_X32 FILLER_17_142 ();
 FILLCELL_X8 FILLER_17_17 ();
 FILLCELL_X8 FILLER_17_174 ();
 FILLCELL_X4 FILLER_17_182 ();
 FILLCELL_X4 FILLER_17_196 ();
 FILLCELL_X1 FILLER_17_200 ();
 FILLCELL_X16 FILLER_17_217 ();
 FILLCELL_X8 FILLER_17_233 ();
 FILLCELL_X4 FILLER_17_241 ();
 FILLCELL_X4 FILLER_17_25 ();
 FILLCELL_X1 FILLER_17_29 ();
 FILLCELL_X32 FILLER_17_46 ();
 FILLCELL_X32 FILLER_17_78 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X1 FILLER_18_103 ();
 FILLCELL_X1 FILLER_18_104 ();
 FILLCELL_X1 FILLER_18_115 ();
 FILLCELL_X1 FILLER_18_116 ();
 FILLCELL_X1 FILLER_18_117 ();
 FILLCELL_X1 FILLER_18_120 ();
 FILLCELL_X1 FILLER_18_121 ();
 FILLCELL_X8 FILLER_18_138 ();
 FILLCELL_X16 FILLER_18_148 ();
 FILLCELL_X4 FILLER_18_164 ();
 FILLCELL_X1 FILLER_18_168 ();
 FILLCELL_X8 FILLER_18_185 ();
 FILLCELL_X1 FILLER_18_193 ();
 FILLCELL_X1 FILLER_18_194 ();
 FILLCELL_X1 FILLER_18_195 ();
 FILLCELL_X32 FILLER_18_198 ();
 FILLCELL_X8 FILLER_18_230 ();
 FILLCELL_X4 FILLER_18_238 ();
 FILLCELL_X1 FILLER_18_242 ();
 FILLCELL_X1 FILLER_18_243 ();
 FILLCELL_X1 FILLER_18_244 ();
 FILLCELL_X16 FILLER_18_33 ();
 FILLCELL_X1 FILLER_18_49 ();
 FILLCELL_X1 FILLER_18_50 ();
 FILLCELL_X16 FILLER_18_53 ();
 FILLCELL_X8 FILLER_18_69 ();
 FILLCELL_X4 FILLER_18_77 ();
 FILLCELL_X1 FILLER_18_81 ();
 FILLCELL_X1 FILLER_18_82 ();
 FILLCELL_X1 FILLER_18_83 ();
 FILLCELL_X8 FILLER_18_87 ();
 FILLCELL_X1 FILLER_18_97 ();
 FILLCELL_X1 FILLER_18_98 ();
 FILLCELL_X1 FILLER_18_99 ();
 FILLCELL_X1 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_100 ();
 FILLCELL_X32 FILLER_19_132 ();
 FILLCELL_X1 FILLER_19_167 ();
 FILLCELL_X1 FILLER_19_168 ();
 FILLCELL_X32 FILLER_19_171 ();
 FILLCELL_X1 FILLER_19_2 ();
 FILLCELL_X32 FILLER_19_203 ();
 FILLCELL_X8 FILLER_19_235 ();
 FILLCELL_X1 FILLER_19_243 ();
 FILLCELL_X1 FILLER_19_244 ();
 FILLCELL_X16 FILLER_19_39 ();
 FILLCELL_X1 FILLER_19_55 ();
 FILLCELL_X1 FILLER_19_56 ();
 FILLCELL_X1 FILLER_19_57 ();
 FILLCELL_X32 FILLER_19_68 ();
 FILLCELL_X32 FILLER_19_7 ();
 FILLCELL_X16 FILLER_1_1 ();
 FILLCELL_X1 FILLER_1_103 ();
 FILLCELL_X1 FILLER_1_104 ();
 FILLCELL_X1 FILLER_1_105 ();
 FILLCELL_X32 FILLER_1_109 ();
 FILLCELL_X32 FILLER_1_141 ();
 FILLCELL_X4 FILLER_1_17 ();
 FILLCELL_X32 FILLER_1_173 ();
 FILLCELL_X16 FILLER_1_205 ();
 FILLCELL_X8 FILLER_1_221 ();
 FILLCELL_X4 FILLER_1_229 ();
 FILLCELL_X1 FILLER_1_233 ();
 FILLCELL_X1 FILLER_1_234 ();
 FILLCELL_X1 FILLER_1_238 ();
 FILLCELL_X1 FILLER_1_239 ();
 FILLCELL_X1 FILLER_1_243 ();
 FILLCELL_X1 FILLER_1_244 ();
 FILLCELL_X32 FILLER_1_25 ();
 FILLCELL_X4 FILLER_1_57 ();
 FILLCELL_X1 FILLER_1_61 ();
 FILLCELL_X32 FILLER_1_67 ();
 FILLCELL_X4 FILLER_1_99 ();
 FILLCELL_X1 FILLER_20_1 ();
 FILLCELL_X1 FILLER_20_112 ();
 FILLCELL_X1 FILLER_20_113 ();
 FILLCELL_X16 FILLER_20_124 ();
 FILLCELL_X4 FILLER_20_140 ();
 FILLCELL_X1 FILLER_20_144 ();
 FILLCELL_X8 FILLER_20_155 ();
 FILLCELL_X4 FILLER_20_163 ();
 FILLCELL_X1 FILLER_20_167 ();
 FILLCELL_X32 FILLER_20_170 ();
 FILLCELL_X1 FILLER_20_2 ();
 FILLCELL_X32 FILLER_20_202 ();
 FILLCELL_X8 FILLER_20_23 ();
 FILLCELL_X8 FILLER_20_234 ();
 FILLCELL_X1 FILLER_20_242 ();
 FILLCELL_X1 FILLER_20_243 ();
 FILLCELL_X1 FILLER_20_244 ();
 FILLCELL_X16 FILLER_20_34 ();
 FILLCELL_X1 FILLER_20_50 ();
 FILLCELL_X1 FILLER_20_51 ();
 FILLCELL_X1 FILLER_20_55 ();
 FILLCELL_X1 FILLER_20_56 ();
 FILLCELL_X8 FILLER_20_59 ();
 FILLCELL_X4 FILLER_20_67 ();
 FILLCELL_X16 FILLER_20_7 ();
 FILLCELL_X1 FILLER_20_71 ();
 FILLCELL_X1 FILLER_20_74 ();
 FILLCELL_X1 FILLER_20_75 ();
 FILLCELL_X8 FILLER_20_79 ();
 FILLCELL_X4 FILLER_20_87 ();
 FILLCELL_X1 FILLER_20_91 ();
 FILLCELL_X1 FILLER_20_92 ();
 FILLCELL_X1 FILLER_20_93 ();
 FILLCELL_X16 FILLER_20_96 ();
 FILLCELL_X1 FILLER_21_1 ();
 FILLCELL_X4 FILLER_21_100 ();
 FILLCELL_X1 FILLER_21_104 ();
 FILLCELL_X1 FILLER_21_105 ();
 FILLCELL_X8 FILLER_21_108 ();
 FILLCELL_X1 FILLER_21_116 ();
 FILLCELL_X1 FILLER_21_117 ();
 FILLCELL_X4 FILLER_21_134 ();
 FILLCELL_X1 FILLER_21_138 ();
 FILLCELL_X1 FILLER_21_139 ();
 FILLCELL_X1 FILLER_21_14 ();
 FILLCELL_X1 FILLER_21_140 ();
 FILLCELL_X1 FILLER_21_15 ();
 FILLCELL_X32 FILLER_21_157 ();
 FILLCELL_X32 FILLER_21_189 ();
 FILLCELL_X1 FILLER_21_2 ();
 FILLCELL_X1 FILLER_21_20 ();
 FILLCELL_X1 FILLER_21_21 ();
 FILLCELL_X16 FILLER_21_221 ();
 FILLCELL_X8 FILLER_21_237 ();
 FILLCELL_X1 FILLER_21_25 ();
 FILLCELL_X1 FILLER_21_26 ();
 FILLCELL_X1 FILLER_21_43 ();
 FILLCELL_X1 FILLER_21_44 ();
 FILLCELL_X16 FILLER_21_47 ();
 FILLCELL_X4 FILLER_21_63 ();
 FILLCELL_X1 FILLER_21_67 ();
 FILLCELL_X1 FILLER_21_68 ();
 FILLCELL_X1 FILLER_21_69 ();
 FILLCELL_X1 FILLER_21_8 ();
 FILLCELL_X1 FILLER_21_86 ();
 FILLCELL_X1 FILLER_21_87 ();
 FILLCELL_X1 FILLER_21_9 ();
 FILLCELL_X4 FILLER_21_90 ();
 FILLCELL_X1 FILLER_21_94 ();
 FILLCELL_X1 FILLER_21_95 ();
 FILLCELL_X1 FILLER_21_96 ();
 FILLCELL_X1 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_109 ();
 FILLCELL_X32 FILLER_22_13 ();
 FILLCELL_X4 FILLER_22_141 ();
 FILLCELL_X1 FILLER_22_145 ();
 FILLCELL_X1 FILLER_22_149 ();
 FILLCELL_X1 FILLER_22_150 ();
 FILLCELL_X32 FILLER_22_153 ();
 FILLCELL_X32 FILLER_22_185 ();
 FILLCELL_X1 FILLER_22_2 ();
 FILLCELL_X16 FILLER_22_217 ();
 FILLCELL_X8 FILLER_22_233 ();
 FILLCELL_X4 FILLER_22_241 ();
 FILLCELL_X32 FILLER_22_45 ();
 FILLCELL_X1 FILLER_22_7 ();
 FILLCELL_X32 FILLER_22_77 ();
 FILLCELL_X1 FILLER_22_8 ();
 FILLCELL_X1 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_103 ();
 FILLCELL_X32 FILLER_23_135 ();
 FILLCELL_X32 FILLER_23_167 ();
 FILLCELL_X32 FILLER_23_199 ();
 FILLCELL_X1 FILLER_23_2 ();
 FILLCELL_X8 FILLER_23_231 ();
 FILLCELL_X4 FILLER_23_239 ();
 FILLCELL_X1 FILLER_23_243 ();
 FILLCELL_X1 FILLER_23_244 ();
 FILLCELL_X32 FILLER_23_39 ();
 FILLCELL_X32 FILLER_23_7 ();
 FILLCELL_X32 FILLER_23_71 ();
 FILLCELL_X16 FILLER_2_1 ();
 FILLCELL_X1 FILLER_2_100 ();
 FILLCELL_X4 FILLER_2_105 ();
 FILLCELL_X1 FILLER_2_109 ();
 FILLCELL_X1 FILLER_2_114 ();
 FILLCELL_X1 FILLER_2_115 ();
 FILLCELL_X8 FILLER_2_119 ();
 FILLCELL_X16 FILLER_2_130 ();
 FILLCELL_X8 FILLER_2_146 ();
 FILLCELL_X1 FILLER_2_154 ();
 FILLCELL_X8 FILLER_2_158 ();
 FILLCELL_X1 FILLER_2_166 ();
 FILLCELL_X1 FILLER_2_167 ();
 FILLCELL_X1 FILLER_2_168 ();
 FILLCELL_X1 FILLER_2_17 ();
 FILLCELL_X1 FILLER_2_171 ();
 FILLCELL_X1 FILLER_2_172 ();
 FILLCELL_X1 FILLER_2_177 ();
 FILLCELL_X1 FILLER_2_178 ();
 FILLCELL_X1 FILLER_2_18 ();
 FILLCELL_X1 FILLER_2_182 ();
 FILLCELL_X1 FILLER_2_183 ();
 FILLCELL_X16 FILLER_2_187 ();
 FILLCELL_X8 FILLER_2_203 ();
 FILLCELL_X4 FILLER_2_211 ();
 FILLCELL_X1 FILLER_2_215 ();
 FILLCELL_X1 FILLER_2_216 ();
 FILLCELL_X1 FILLER_2_217 ();
 FILLCELL_X1 FILLER_2_221 ();
 FILLCELL_X1 FILLER_2_222 ();
 FILLCELL_X1 FILLER_2_226 ();
 FILLCELL_X1 FILLER_2_227 ();
 FILLCELL_X4 FILLER_2_231 ();
 FILLCELL_X1 FILLER_2_238 ();
 FILLCELL_X1 FILLER_2_239 ();
 FILLCELL_X1 FILLER_2_243 ();
 FILLCELL_X1 FILLER_2_244 ();
 FILLCELL_X1 FILLER_2_28 ();
 FILLCELL_X1 FILLER_2_29 ();
 FILLCELL_X4 FILLER_2_32 ();
 FILLCELL_X1 FILLER_2_36 ();
 FILLCELL_X1 FILLER_2_37 ();
 FILLCELL_X8 FILLER_2_41 ();
 FILLCELL_X4 FILLER_2_49 ();
 FILLCELL_X1 FILLER_2_62 ();
 FILLCELL_X1 FILLER_2_63 ();
 FILLCELL_X1 FILLER_2_73 ();
 FILLCELL_X1 FILLER_2_74 ();
 FILLCELL_X16 FILLER_2_79 ();
 FILLCELL_X4 FILLER_2_95 ();
 FILLCELL_X1 FILLER_2_99 ();
 FILLCELL_X16 FILLER_3_1 ();
 FILLCELL_X1 FILLER_3_102 ();
 FILLCELL_X1 FILLER_3_103 ();
 FILLCELL_X1 FILLER_3_104 ();
 FILLCELL_X1 FILLER_3_109 ();
 FILLCELL_X1 FILLER_3_110 ();
 FILLCELL_X1 FILLER_3_114 ();
 FILLCELL_X1 FILLER_3_115 ();
 FILLCELL_X16 FILLER_3_119 ();
 FILLCELL_X8 FILLER_3_135 ();
 FILLCELL_X4 FILLER_3_143 ();
 FILLCELL_X1 FILLER_3_147 ();
 FILLCELL_X1 FILLER_3_148 ();
 FILLCELL_X4 FILLER_3_153 ();
 FILLCELL_X1 FILLER_3_161 ();
 FILLCELL_X1 FILLER_3_162 ();
 FILLCELL_X1 FILLER_3_166 ();
 FILLCELL_X1 FILLER_3_167 ();
 FILLCELL_X8 FILLER_3_17 ();
 FILLCELL_X1 FILLER_3_170 ();
 FILLCELL_X1 FILLER_3_171 ();
 FILLCELL_X1 FILLER_3_174 ();
 FILLCELL_X1 FILLER_3_175 ();
 FILLCELL_X1 FILLER_3_180 ();
 FILLCELL_X1 FILLER_3_181 ();
 FILLCELL_X1 FILLER_3_186 ();
 FILLCELL_X1 FILLER_3_187 ();
 FILLCELL_X16 FILLER_3_192 ();
 FILLCELL_X8 FILLER_3_208 ();
 FILLCELL_X1 FILLER_3_218 ();
 FILLCELL_X1 FILLER_3_219 ();
 FILLCELL_X1 FILLER_3_220 ();
 FILLCELL_X16 FILLER_3_223 ();
 FILLCELL_X1 FILLER_3_239 ();
 FILLCELL_X1 FILLER_3_243 ();
 FILLCELL_X1 FILLER_3_244 ();
 FILLCELL_X4 FILLER_3_25 ();
 FILLCELL_X4 FILLER_3_32 ();
 FILLCELL_X1 FILLER_3_36 ();
 FILLCELL_X1 FILLER_3_37 ();
 FILLCELL_X1 FILLER_3_38 ();
 FILLCELL_X16 FILLER_3_44 ();
 FILLCELL_X8 FILLER_3_60 ();
 FILLCELL_X1 FILLER_3_68 ();
 FILLCELL_X16 FILLER_3_73 ();
 FILLCELL_X4 FILLER_3_89 ();
 FILLCELL_X1 FILLER_3_95 ();
 FILLCELL_X1 FILLER_3_96 ();
 FILLCELL_X1 FILLER_3_97 ();
 FILLCELL_X8 FILLER_4_1 ();
 FILLCELL_X1 FILLER_4_10 ();
 FILLCELL_X1 FILLER_4_11 ();
 FILLCELL_X8 FILLER_4_131 ();
 FILLCELL_X1 FILLER_4_139 ();
 FILLCELL_X1 FILLER_4_140 ();
 FILLCELL_X1 FILLER_4_145 ();
 FILLCELL_X1 FILLER_4_146 ();
 FILLCELL_X1 FILLER_4_150 ();
 FILLCELL_X1 FILLER_4_151 ();
 FILLCELL_X8 FILLER_4_154 ();
 FILLCELL_X4 FILLER_4_162 ();
 FILLCELL_X1 FILLER_4_166 ();
 FILLCELL_X1 FILLER_4_167 ();
 FILLCELL_X1 FILLER_4_17 ();
 FILLCELL_X8 FILLER_4_172 ();
 FILLCELL_X1 FILLER_4_18 ();
 FILLCELL_X1 FILLER_4_180 ();
 FILLCELL_X32 FILLER_4_184 ();
 FILLCELL_X16 FILLER_4_216 ();
 FILLCELL_X8 FILLER_4_232 ();
 FILLCELL_X4 FILLER_4_240 ();
 FILLCELL_X1 FILLER_4_244 ();
 FILLCELL_X1 FILLER_4_28 ();
 FILLCELL_X1 FILLER_4_29 ();
 FILLCELL_X1 FILLER_4_35 ();
 FILLCELL_X1 FILLER_4_36 ();
 FILLCELL_X32 FILLER_4_40 ();
 FILLCELL_X16 FILLER_4_72 ();
 FILLCELL_X4 FILLER_4_88 ();
 FILLCELL_X1 FILLER_4_9 ();
 FILLCELL_X1 FILLER_4_92 ();
 FILLCELL_X1 FILLER_4_93 ();
 FILLCELL_X1 FILLER_4_94 ();
 FILLCELL_X32 FILLER_4_99 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_112 ();
 FILLCELL_X4 FILLER_5_144 ();
 FILLCELL_X1 FILLER_5_148 ();
 FILLCELL_X32 FILLER_5_159 ();
 FILLCELL_X32 FILLER_5_191 ();
 FILLCELL_X16 FILLER_5_223 ();
 FILLCELL_X4 FILLER_5_239 ();
 FILLCELL_X1 FILLER_5_243 ();
 FILLCELL_X1 FILLER_5_244 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X8 FILLER_5_65 ();
 FILLCELL_X1 FILLER_5_73 ();
 FILLCELL_X1 FILLER_5_74 ();
 FILLCELL_X1 FILLER_5_75 ();
 FILLCELL_X32 FILLER_5_80 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_102 ();
 FILLCELL_X32 FILLER_6_134 ();
 FILLCELL_X32 FILLER_6_166 ();
 FILLCELL_X32 FILLER_6_198 ();
 FILLCELL_X8 FILLER_6_230 ();
 FILLCELL_X4 FILLER_6_238 ();
 FILLCELL_X1 FILLER_6_242 ();
 FILLCELL_X1 FILLER_6_243 ();
 FILLCELL_X1 FILLER_6_244 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X1 FILLER_6_97 ();
 FILLCELL_X1 FILLER_6_98 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X1 FILLER_7_102 ();
 FILLCELL_X1 FILLER_7_103 ();
 FILLCELL_X32 FILLER_7_108 ();
 FILLCELL_X32 FILLER_7_140 ();
 FILLCELL_X16 FILLER_7_172 ();
 FILLCELL_X1 FILLER_7_188 ();
 FILLCELL_X1 FILLER_7_189 ();
 FILLCELL_X1 FILLER_7_190 ();
 FILLCELL_X1 FILLER_7_193 ();
 FILLCELL_X1 FILLER_7_194 ();
 FILLCELL_X1 FILLER_7_199 ();
 FILLCELL_X1 FILLER_7_200 ();
 FILLCELL_X1 FILLER_7_204 ();
 FILLCELL_X1 FILLER_7_205 ();
 FILLCELL_X1 FILLER_7_209 ();
 FILLCELL_X1 FILLER_7_210 ();
 FILLCELL_X8 FILLER_7_214 ();
 FILLCELL_X16 FILLER_7_226 ();
 FILLCELL_X1 FILLER_7_242 ();
 FILLCELL_X1 FILLER_7_243 ();
 FILLCELL_X1 FILLER_7_244 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X16 FILLER_7_65 ();
 FILLCELL_X1 FILLER_7_81 ();
 FILLCELL_X1 FILLER_7_82 ();
 FILLCELL_X1 FILLER_7_83 ();
 FILLCELL_X4 FILLER_7_94 ();
 FILLCELL_X16 FILLER_8_1 ();
 FILLCELL_X8 FILLER_8_122 ();
 FILLCELL_X1 FILLER_8_130 ();
 FILLCELL_X8 FILLER_8_135 ();
 FILLCELL_X4 FILLER_8_143 ();
 FILLCELL_X1 FILLER_8_147 ();
 FILLCELL_X1 FILLER_8_148 ();
 FILLCELL_X32 FILLER_8_153 ();
 FILLCELL_X8 FILLER_8_17 ();
 FILLCELL_X1 FILLER_8_185 ();
 FILLCELL_X1 FILLER_8_186 ();
 FILLCELL_X1 FILLER_8_191 ();
 FILLCELL_X1 FILLER_8_192 ();
 FILLCELL_X1 FILLER_8_193 ();
 FILLCELL_X1 FILLER_8_198 ();
 FILLCELL_X1 FILLER_8_199 ();
 FILLCELL_X1 FILLER_8_204 ();
 FILLCELL_X1 FILLER_8_205 ();
 FILLCELL_X1 FILLER_8_210 ();
 FILLCELL_X1 FILLER_8_211 ();
 FILLCELL_X16 FILLER_8_215 ();
 FILLCELL_X8 FILLER_8_231 ();
 FILLCELL_X1 FILLER_8_239 ();
 FILLCELL_X1 FILLER_8_243 ();
 FILLCELL_X1 FILLER_8_244 ();
 FILLCELL_X1 FILLER_8_25 ();
 FILLCELL_X8 FILLER_8_28 ();
 FILLCELL_X1 FILLER_8_39 ();
 FILLCELL_X1 FILLER_8_40 ();
 FILLCELL_X1 FILLER_8_44 ();
 FILLCELL_X1 FILLER_8_45 ();
 FILLCELL_X1 FILLER_8_46 ();
 FILLCELL_X4 FILLER_8_49 ();
 FILLCELL_X1 FILLER_8_53 ();
 FILLCELL_X32 FILLER_8_58 ();
 FILLCELL_X32 FILLER_8_90 ();
 FILLCELL_X16 FILLER_9_1 ();
 FILLCELL_X1 FILLER_9_100 ();
 FILLCELL_X16 FILLER_9_103 ();
 FILLCELL_X4 FILLER_9_119 ();
 FILLCELL_X1 FILLER_9_123 ();
 FILLCELL_X1 FILLER_9_124 ();
 FILLCELL_X1 FILLER_9_125 ();
 FILLCELL_X16 FILLER_9_130 ();
 FILLCELL_X1 FILLER_9_146 ();
 FILLCELL_X1 FILLER_9_147 ();
 FILLCELL_X8 FILLER_9_151 ();
 FILLCELL_X1 FILLER_9_159 ();
 FILLCELL_X16 FILLER_9_162 ();
 FILLCELL_X4 FILLER_9_17 ();
 FILLCELL_X4 FILLER_9_178 ();
 FILLCELL_X1 FILLER_9_182 ();
 FILLCELL_X1 FILLER_9_183 ();
 FILLCELL_X1 FILLER_9_188 ();
 FILLCELL_X1 FILLER_9_189 ();
 FILLCELL_X1 FILLER_9_200 ();
 FILLCELL_X1 FILLER_9_201 ();
 FILLCELL_X16 FILLER_9_205 ();
 FILLCELL_X1 FILLER_9_221 ();
 FILLCELL_X1 FILLER_9_222 ();
 FILLCELL_X8 FILLER_9_225 ();
 FILLCELL_X4 FILLER_9_233 ();
 FILLCELL_X1 FILLER_9_237 ();
 FILLCELL_X1 FILLER_9_238 ();
 FILLCELL_X1 FILLER_9_239 ();
 FILLCELL_X1 FILLER_9_24 ();
 FILLCELL_X1 FILLER_9_243 ();
 FILLCELL_X1 FILLER_9_244 ();
 FILLCELL_X1 FILLER_9_25 ();
 FILLCELL_X4 FILLER_9_30 ();
 FILLCELL_X1 FILLER_9_34 ();
 FILLCELL_X1 FILLER_9_39 ();
 FILLCELL_X1 FILLER_9_40 ();
 FILLCELL_X1 FILLER_9_41 ();
 FILLCELL_X4 FILLER_9_46 ();
 FILLCELL_X1 FILLER_9_50 ();
 FILLCELL_X1 FILLER_9_55 ();
 FILLCELL_X1 FILLER_9_56 ();
 FILLCELL_X1 FILLER_9_60 ();
 FILLCELL_X1 FILLER_9_61 ();
 FILLCELL_X16 FILLER_9_65 ();
 FILLCELL_X4 FILLER_9_81 ();
 FILLCELL_X1 FILLER_9_85 ();
 FILLCELL_X1 FILLER_9_86 ();
 FILLCELL_X8 FILLER_9_91 ();
 FILLCELL_X1 FILLER_9_99 ();
 TAPCELL_X1 PHY_0 ();
 TAPCELL_X1 PHY_1 ();
 TAPCELL_X1 PHY_10 ();
 TAPCELL_X1 PHY_11 ();
 TAPCELL_X1 PHY_12 ();
 TAPCELL_X1 PHY_13 ();
 TAPCELL_X1 PHY_14 ();
 TAPCELL_X1 PHY_15 ();
 TAPCELL_X1 PHY_16 ();
 TAPCELL_X1 PHY_17 ();
 TAPCELL_X1 PHY_18 ();
 TAPCELL_X1 PHY_19 ();
 TAPCELL_X1 PHY_2 ();
 TAPCELL_X1 PHY_20 ();
 TAPCELL_X1 PHY_21 ();
 TAPCELL_X1 PHY_22 ();
 TAPCELL_X1 PHY_23 ();
 TAPCELL_X1 PHY_24 ();
 TAPCELL_X1 PHY_25 ();
 TAPCELL_X1 PHY_26 ();
 TAPCELL_X1 PHY_27 ();
 TAPCELL_X1 PHY_28 ();
 TAPCELL_X1 PHY_29 ();
 TAPCELL_X1 PHY_3 ();
 TAPCELL_X1 PHY_30 ();
 TAPCELL_X1 PHY_31 ();
 TAPCELL_X1 PHY_32 ();
 TAPCELL_X1 PHY_33 ();
 TAPCELL_X1 PHY_34 ();
 TAPCELL_X1 PHY_35 ();
 TAPCELL_X1 PHY_36 ();
 TAPCELL_X1 PHY_37 ();
 TAPCELL_X1 PHY_38 ();
 TAPCELL_X1 PHY_39 ();
 TAPCELL_X1 PHY_4 ();
 TAPCELL_X1 PHY_40 ();
 TAPCELL_X1 PHY_41 ();
 TAPCELL_X1 PHY_42 ();
 TAPCELL_X1 PHY_43 ();
 TAPCELL_X1 PHY_44 ();
 TAPCELL_X1 PHY_45 ();
 TAPCELL_X1 PHY_46 ();
 TAPCELL_X1 PHY_47 ();
 TAPCELL_X1 PHY_5 ();
 TAPCELL_X1 PHY_6 ();
 TAPCELL_X1 PHY_7 ();
 TAPCELL_X1 PHY_8 ();
 TAPCELL_X1 PHY_9 ();
 INV_X4 _201_ (.A(net11),
    .ZN(_107_));
 NOR2_X4 _203_ (.A1(_107_),
    .A2(net12),
    .ZN(_109_));
 INV_X2 _206_ (.A(net10),
    .ZN(_112_));
 NOR2_X2 _208_ (.A1(_112_),
    .A2(net9),
    .ZN(_001_));
 NAND3_X1 _209_ (.A1(_109_),
    .A2(_001_),
    .A3(_171_),
    .ZN(_002_));
 NAND2_X1 _210_ (.A1(net9),
    .A2(net10),
    .ZN(_003_));
 INV_X2 _211_ (.A(_003_),
    .ZN(_004_));
 NOR2_X4 _212_ (.A1(net11),
    .A2(net12),
    .ZN(_005_));
 NAND2_X1 _213_ (.A1(_004_),
    .A2(_005_),
    .ZN(_006_));
 OAI21_X1 _214_ (.A(_002_),
    .B1(_171_),
    .B2(_006_),
    .ZN(_007_));
 INV_X4 _215_ (.A(net9),
    .ZN(_008_));
 NOR2_X4 _216_ (.A1(_008_),
    .A2(net10),
    .ZN(_009_));
 INV_X1 _217_ (.A(_162_),
    .ZN(_010_));
 NAND3_X1 _218_ (.A1(_009_),
    .A2(_109_),
    .A3(_010_),
    .ZN(_011_));
 NAND3_X1 _219_ (.A1(_109_),
    .A2(_004_),
    .A3(_172_),
    .ZN(_012_));
 INV_X1 _220_ (.A(net12),
    .ZN(_013_));
 NOR2_X4 _221_ (.A1(_013_),
    .A2(net11),
    .ZN(_014_));
 NOR2_X2 _222_ (.A1(net9),
    .A2(net10),
    .ZN(_015_));
 INV_X1 _223_ (.A(_172_),
    .ZN(_016_));
 NAND3_X1 _224_ (.A1(_014_),
    .A2(_015_),
    .A3(_016_),
    .ZN(_017_));
 NAND3_X1 _225_ (.A1(_011_),
    .A2(_012_),
    .A3(_017_),
    .ZN(_018_));
 NOR2_X1 _226_ (.A1(_007_),
    .A2(_018_),
    .ZN(_019_));
 INV_X1 _227_ (.A(net1),
    .ZN(_169_));
 NAND3_X1 _228_ (.A1(_109_),
    .A2(_015_),
    .A3(_169_),
    .ZN(_020_));
 NAND3_X1 _229_ (.A1(_112_),
    .A2(_107_),
    .A3(_172_),
    .ZN(_021_));
 OAI21_X1 _230_ (.A(_020_),
    .B1(net12),
    .B2(_021_),
    .ZN(_022_));
 NAND2_X1 _231_ (.A1(_009_),
    .A2(_014_),
    .ZN(_023_));
 NAND2_X1 _232_ (.A1(_001_),
    .A2(_005_),
    .ZN(_024_));
 AOI21_X1 _233_ (.A(_010_),
    .B1(_023_),
    .B2(_024_),
    .ZN(_025_));
 NOR2_X1 _234_ (.A1(_022_),
    .A2(_025_),
    .ZN(_026_));
 NAND2_X1 _235_ (.A1(_019_),
    .A2(_026_),
    .ZN(net13));
 NAND2_X1 _236_ (.A1(net2),
    .A2(net5),
    .ZN(_027_));
 INV_X1 _237_ (.A(_027_),
    .ZN(_177_));
 INV_X1 _238_ (.A(_183_),
    .ZN(_167_));
 NAND3_X1 _239_ (.A1(_109_),
    .A2(_001_),
    .A3(_181_),
    .ZN(_028_));
 NAND3_X1 _240_ (.A1(_109_),
    .A2(_004_),
    .A3(_182_),
    .ZN(_029_));
 NAND2_X1 _241_ (.A1(_028_),
    .A2(_029_),
    .ZN(_030_));
 NAND3_X1 _242_ (.A1(_009_),
    .A2(_014_),
    .A3(_179_),
    .ZN(_031_));
 INV_X1 _243_ (.A(_182_),
    .ZN(_032_));
 NAND3_X1 _244_ (.A1(_014_),
    .A2(_015_),
    .A3(_032_),
    .ZN(_033_));
 NAND2_X1 _245_ (.A1(_031_),
    .A2(_033_),
    .ZN(_034_));
 NOR2_X1 _246_ (.A1(_030_),
    .A2(_034_),
    .ZN(_035_));
 NAND3_X1 _247_ (.A1(_009_),
    .A2(_109_),
    .A3(_167_),
    .ZN(_036_));
 INV_X1 _248_ (.A(net2),
    .ZN(_180_));
 NAND3_X1 _249_ (.A1(_109_),
    .A2(_015_),
    .A3(_180_),
    .ZN(_037_));
 NAND2_X1 _250_ (.A1(_036_),
    .A2(_037_),
    .ZN(_038_));
 INV_X1 _251_ (.A(_181_),
    .ZN(_039_));
 NAND3_X1 _252_ (.A1(_004_),
    .A2(_005_),
    .A3(_039_),
    .ZN(_040_));
 NAND3_X1 _253_ (.A1(_001_),
    .A2(_005_),
    .A3(_183_),
    .ZN(_041_));
 NAND2_X1 _254_ (.A1(_040_),
    .A2(_041_),
    .ZN(_042_));
 NOR2_X1 _255_ (.A1(_038_),
    .A2(_042_),
    .ZN(_043_));
 AND2_X1 _256_ (.A1(_009_),
    .A2(_005_),
    .ZN(_044_));
 NAND2_X1 _257_ (.A1(_044_),
    .A2(_161_),
    .ZN(_045_));
 AND2_X1 _258_ (.A1(_005_),
    .A2(_015_),
    .ZN(_046_));
 NAND2_X1 _259_ (.A1(_046_),
    .A2(_164_),
    .ZN(_047_));
 NAND2_X1 _260_ (.A1(_045_),
    .A2(_047_),
    .ZN(_048_));
 INV_X1 _261_ (.A(_048_),
    .ZN(_049_));
 NAND3_X1 _262_ (.A1(_035_),
    .A2(_043_),
    .A3(_049_),
    .ZN(net14));
 NAND3_X1 _263_ (.A1(_109_),
    .A2(_001_),
    .A3(_189_),
    .ZN(_050_));
 NAND3_X1 _264_ (.A1(_109_),
    .A2(_004_),
    .A3(_190_),
    .ZN(_051_));
 NAND2_X1 _265_ (.A1(_050_),
    .A2(_051_),
    .ZN(_052_));
 NAND3_X1 _266_ (.A1(_009_),
    .A2(_014_),
    .A3(_188_),
    .ZN(_053_));
 INV_X1 _267_ (.A(_190_),
    .ZN(_054_));
 NAND3_X1 _268_ (.A1(_014_),
    .A2(_015_),
    .A3(_054_),
    .ZN(_055_));
 NAND2_X1 _269_ (.A1(_053_),
    .A2(_055_),
    .ZN(_056_));
 NOR2_X1 _270_ (.A1(_052_),
    .A2(_056_),
    .ZN(_057_));
 INV_X1 _271_ (.A(_138_),
    .ZN(_058_));
 NAND3_X1 _272_ (.A1(_009_),
    .A2(_109_),
    .A3(_058_),
    .ZN(_059_));
 INV_X1 _273_ (.A(net3),
    .ZN(_117_));
 NAND3_X1 _274_ (.A1(_109_),
    .A2(_015_),
    .A3(_117_),
    .ZN(_060_));
 NAND2_X1 _275_ (.A1(_059_),
    .A2(_060_),
    .ZN(_061_));
 NAND3_X1 _276_ (.A1(_001_),
    .A2(_005_),
    .A3(_138_),
    .ZN(_062_));
 INV_X1 _277_ (.A(_189_),
    .ZN(_063_));
 NAND3_X1 _278_ (.A1(_004_),
    .A2(_005_),
    .A3(_063_),
    .ZN(_064_));
 NAND2_X1 _279_ (.A1(_062_),
    .A2(_064_),
    .ZN(_065_));
 NOR2_X1 _280_ (.A1(_061_),
    .A2(_065_),
    .ZN(_066_));
 NAND2_X1 _281_ (.A1(_044_),
    .A2(_116_),
    .ZN(_067_));
 INV_X1 _282_ (.A(_120_),
    .ZN(_068_));
 NAND2_X1 _283_ (.A1(_046_),
    .A2(_068_),
    .ZN(_069_));
 NAND2_X1 _284_ (.A1(_067_),
    .A2(_069_),
    .ZN(_070_));
 INV_X1 _285_ (.A(_070_),
    .ZN(_071_));
 NAND3_X1 _286_ (.A1(_057_),
    .A2(_066_),
    .A3(_071_),
    .ZN(net15));
 NAND2_X1 _287_ (.A1(net1),
    .A2(net8),
    .ZN(_072_));
 INV_X1 _288_ (.A(_072_),
    .ZN(_192_));
 NAND2_X1 _289_ (.A1(net2),
    .A2(net7),
    .ZN(_127_));
 NAND2_X1 _290_ (.A1(net5),
    .A2(net4),
    .ZN(_121_));
 NAND2_X1 _291_ (.A1(net6),
    .A2(net3),
    .ZN(_123_));
 NAND3_X1 _292_ (.A1(_109_),
    .A2(_001_),
    .A3(_195_),
    .ZN(_073_));
 NAND3_X1 _293_ (.A1(_109_),
    .A2(_004_),
    .A3(_196_),
    .ZN(_074_));
 NAND2_X1 _294_ (.A1(_073_),
    .A2(_074_),
    .ZN(_075_));
 NAND3_X1 _295_ (.A1(_009_),
    .A2(_014_),
    .A3(_194_),
    .ZN(_076_));
 INV_X1 _296_ (.A(_196_),
    .ZN(_077_));
 NAND3_X1 _297_ (.A1(_014_),
    .A2(_015_),
    .A3(_077_),
    .ZN(_078_));
 NAND2_X1 _298_ (.A1(_076_),
    .A2(_078_),
    .ZN(_079_));
 NOR2_X1 _299_ (.A1(_075_),
    .A2(_079_),
    .ZN(_080_));
 INV_X1 _300_ (.A(_156_),
    .ZN(_081_));
 NAND3_X1 _301_ (.A1(_009_),
    .A2(_109_),
    .A3(_081_),
    .ZN(_082_));
 INV_X2 _302_ (.A(net4),
    .ZN(_130_));
 NAND3_X1 _303_ (.A1(_109_),
    .A2(_015_),
    .A3(_130_),
    .ZN(_083_));
 NAND2_X1 _304_ (.A1(_082_),
    .A2(_083_),
    .ZN(_084_));
 NAND3_X1 _305_ (.A1(_001_),
    .A2(_005_),
    .A3(_156_),
    .ZN(_085_));
 INV_X1 _306_ (.A(_195_),
    .ZN(_086_));
 NAND3_X1 _307_ (.A1(_004_),
    .A2(_005_),
    .A3(_086_),
    .ZN(_087_));
 NAND2_X1 _308_ (.A1(_085_),
    .A2(_087_),
    .ZN(_088_));
 NOR2_X1 _309_ (.A1(_084_),
    .A2(_088_),
    .ZN(_089_));
 NAND2_X1 _310_ (.A1(_044_),
    .A2(_133_),
    .ZN(_090_));
 INV_X1 _311_ (.A(_136_),
    .ZN(_091_));
 NAND2_X1 _312_ (.A1(_046_),
    .A2(_091_),
    .ZN(_092_));
 NAND2_X1 _313_ (.A1(_090_),
    .A2(_092_),
    .ZN(_093_));
 INV_X1 _314_ (.A(_093_),
    .ZN(_094_));
 NAND3_X1 _315_ (.A1(_080_),
    .A2(_089_),
    .A3(_094_),
    .ZN(net16));
 NAND2_X1 _316_ (.A1(net2),
    .A2(net8),
    .ZN(_095_));
 INV_X1 _317_ (.A(_095_),
    .ZN(_142_));
 NAND2_X1 _318_ (.A1(net6),
    .A2(net4),
    .ZN(_096_));
 INV_X1 _319_ (.A(_096_),
    .ZN(_198_));
 NAND2_X1 _320_ (.A1(_044_),
    .A2(_132_),
    .ZN(_097_));
 INV_X1 _321_ (.A(_135_),
    .ZN(_098_));
 NAND2_X1 _322_ (.A1(_046_),
    .A2(_098_),
    .ZN(_099_));
 NAND3_X1 _323_ (.A1(_009_),
    .A2(_014_),
    .A3(_145_),
    .ZN(_100_));
 NAND3_X1 _324_ (.A1(_097_),
    .A2(_099_),
    .A3(_100_),
    .ZN(net17));
 NAND2_X1 _325_ (.A1(net3),
    .A2(net8),
    .ZN(_152_));
 NAND2_X1 _326_ (.A1(net7),
    .A2(net4),
    .ZN(_101_));
 INV_X1 _327_ (.A(_101_),
    .ZN(_146_));
 NOR2_X1 _328_ (.A1(_023_),
    .A2(_154_),
    .ZN(net18));
 INV_X1 _329_ (.A(_158_),
    .ZN(_102_));
 NOR2_X1 _330_ (.A1(_023_),
    .A2(_102_),
    .ZN(net19));
 INV_X1 _331_ (.A(_157_),
    .ZN(_103_));
 NOR2_X1 _332_ (.A1(_023_),
    .A2(_103_),
    .ZN(net20));
 INV_X1 _333_ (.A(_153_),
    .ZN(_155_));
 NAND2_X1 _334_ (.A1(net5),
    .A2(net3),
    .ZN(_166_));
 INV_X1 _335_ (.A(_149_),
    .ZN(_151_));
 INV_X1 _336_ (.A(_115_),
    .ZN(_131_));
 INV_X1 _337_ (.A(_144_),
    .ZN(_150_));
 INV_X1 _338_ (.A(_163_),
    .ZN(_118_));
 NAND2_X1 _339_ (.A1(net1),
    .A2(net6),
    .ZN(_104_));
 INV_X1 _340_ (.A(_104_),
    .ZN(_176_));
 INV_X1 _341_ (.A(_173_),
    .ZN(_160_));
 NAND2_X1 _342_ (.A1(net1),
    .A2(net7),
    .ZN(_105_));
 INV_X1 _343_ (.A(_105_),
    .ZN(_185_));
 INV_X1 _344_ (.A(net5),
    .ZN(_170_));
 INV_X1 _345_ (.A(net6),
    .ZN(_159_));
 INV_X1 _346_ (.A(_168_),
    .ZN(_186_));
 INV_X1 _347_ (.A(net7),
    .ZN(_113_));
 INV_X1 _348_ (.A(_129_),
    .ZN(_193_));
 INV_X1 _349_ (.A(net8),
    .ZN(_134_));
 INV_X1 _350_ (.A(_124_),
    .ZN(_199_));
 INV_X1 _351_ (.A(_128_),
    .ZN(_139_));
 INV_X1 _352_ (.A(_178_),
    .ZN(_165_));
 INV_X1 _353_ (.A(_187_),
    .ZN(_126_));
 FA_X1 _354_ (.A(net3),
    .B(_113_),
    .CI(_114_),
    .CO(_115_),
    .S(_116_));
 FA_X1 _355_ (.A(_117_),
    .B(_113_),
    .CI(_118_),
    .CO(_119_),
    .S(_120_));
 FA_X1 _356_ (.A(_121_),
    .B(_122_),
    .CI(_123_),
    .CO(_124_),
    .S(_125_));
 FA_X1 _357_ (.A(_126_),
    .B(_125_),
    .CI(_127_),
    .CO(_128_),
    .S(_129_));
 FA_X1 _358_ (.A(_130_),
    .B(net8),
    .CI(_131_),
    .CO(_132_),
    .S(_133_));
 FA_X1 _359_ (.A(_130_),
    .B(_134_),
    .CI(_119_),
    .CO(_135_),
    .S(_136_));
 FA_X1 _360_ (.A(_137_),
    .B(_138_),
    .CI(_139_),
    .CO(_140_),
    .S(_141_));
 FA_X1 _361_ (.A(_141_),
    .B(_142_),
    .CI(_143_),
    .CO(_144_),
    .S(_145_));
 FA_X1 _362_ (.A(_146_),
    .B(_147_),
    .CI(_140_),
    .CO(_148_),
    .S(_149_));
 FA_X1 _363_ (.A(_150_),
    .B(_151_),
    .CI(_152_),
    .CO(_153_),
    .S(_154_));
 FA_X1 _364_ (.A(_155_),
    .B(_148_),
    .CI(_156_),
    .CO(_157_),
    .S(_158_));
 FA_X1 _365_ (.A(net2),
    .B(_159_),
    .CI(_160_),
    .CO(_114_),
    .S(_161_));
 FA_X1 _366_ (.A(net2),
    .B(net6),
    .CI(_162_),
    .CO(_163_),
    .S(_164_));
 FA_X1 _367_ (.A(_165_),
    .B(_166_),
    .CI(_167_),
    .CO(_122_),
    .S(_168_));
 HA_X1 _368_ (.A(_169_),
    .B(_170_),
    .CO(_171_),
    .S(_172_));
 HA_X1 _369_ (.A(_169_),
    .B(net5),
    .CO(_173_),
    .S(_174_));
 HA_X1 _370_ (.A(net1),
    .B(net5),
    .CO(_162_),
    .S(_175_));
 HA_X1 _371_ (.A(_176_),
    .B(_177_),
    .CO(_178_),
    .S(_179_));
 HA_X1 _372_ (.A(_180_),
    .B(_159_),
    .CO(_181_),
    .S(_182_));
 HA_X1 _373_ (.A(net2),
    .B(net6),
    .CO(_183_),
    .S(_184_));
 HA_X1 _374_ (.A(_185_),
    .B(_186_),
    .CO(_187_),
    .S(_188_));
 HA_X1 _375_ (.A(_117_),
    .B(_113_),
    .CO(_189_),
    .S(_190_));
 HA_X1 _376_ (.A(net3),
    .B(net7),
    .CO(_138_),
    .S(_191_));
 HA_X1 _377_ (.A(_192_),
    .B(_193_),
    .CO(_143_),
    .S(_194_));
 HA_X1 _378_ (.A(_130_),
    .B(_134_),
    .CO(_195_),
    .S(_196_));
 HA_X1 _379_ (.A(net4),
    .B(net8),
    .CO(_156_),
    .S(_197_));
 HA_X1 _380_ (.A(_198_),
    .B(_199_),
    .CO(_147_),
    .S(_137_));
 CLKBUF_X2 input1 (.A(A[0]),
    .Z(net1));
 BUF_X2 input10 (.A(CTRL[1]),
    .Z(net10));
 CLKBUF_X3 input11 (.A(CTRL[2]),
    .Z(net11));
 BUF_X2 input12 (.A(CTRL[3]),
    .Z(net12));
 CLKBUF_X3 input2 (.A(A[1]),
    .Z(net2));
 BUF_X2 input3 (.A(A[2]),
    .Z(net3));
 BUF_X2 input4 (.A(A[3]),
    .Z(net4));
 BUF_X2 input5 (.A(B[0]),
    .Z(net5));
 BUF_X2 input6 (.A(B[1]),
    .Z(net6));
 CLKBUF_X2 input7 (.A(B[2]),
    .Z(net7));
 BUF_X2 input8 (.A(B[3]),
    .Z(net8));
 BUF_X2 input9 (.A(CTRL[0]),
    .Z(net9));
 BUF_X1 output13 (.A(net13),
    .Z(Y[0]));
 BUF_X1 output14 (.A(net14),
    .Z(Y[1]));
 BUF_X1 output15 (.A(net15),
    .Z(Y[2]));
 BUF_X1 output16 (.A(net16),
    .Z(Y[3]));
 BUF_X1 output17 (.A(net17),
    .Z(Y[4]));
 BUF_X1 output18 (.A(net18),
    .Z(Y[5]));
 BUF_X1 output19 (.A(net19),
    .Z(Y[6]));
 BUF_X1 output20 (.A(net20),
    .Z(Y[7]));
endmodule

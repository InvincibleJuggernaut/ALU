module alu_4 (A,
    B,
    CTRL,
    Y);
 input [3:0] A;
 input [3:0] B;
 input [3:0] CTRL;
 output [7:0] Y;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _130_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;

 INV_X4 _225_ (.A(CTRL[1]),
    .ZN(_130_));
 NAND2_X1 _227_ (.A1(_130_),
    .A2(CTRL[0]),
    .ZN(_132_));
 INV_X2 _228_ (.A(CTRL[3]),
    .ZN(_000_));
 NAND2_X2 _229_ (.A1(_000_),
    .A2(CTRL[2]),
    .ZN(_001_));
 NOR2_X2 _230_ (.A1(_132_),
    .A2(_001_),
    .ZN(_002_));
 INV_X1 _231_ (.A(_163_),
    .ZN(_003_));
 NAND2_X1 _232_ (.A1(_002_),
    .A2(_003_),
    .ZN(_004_));
 INV_X4 _233_ (.A(CTRL[0]),
    .ZN(_005_));
 NAND2_X1 _234_ (.A1(_005_),
    .A2(CTRL[1]),
    .ZN(_006_));
 NOR2_X2 _235_ (.A1(_006_),
    .A2(_001_),
    .ZN(_007_));
 NAND2_X1 _236_ (.A1(_007_),
    .A2(_206_),
    .ZN(_008_));
 NAND2_X1 _237_ (.A1(_004_),
    .A2(_008_),
    .ZN(_009_));
 NAND2_X1 _238_ (.A1(_130_),
    .A2(_005_),
    .ZN(_010_));
 NOR2_X2 _239_ (.A1(_010_),
    .A2(_001_),
    .ZN(_011_));
 INV_X1 _240_ (.A(A[2]),
    .ZN(_142_));
 NAND2_X1 _241_ (.A1(_011_),
    .A2(_142_),
    .ZN(_012_));
 INV_X2 _242_ (.A(CTRL[2]),
    .ZN(_013_));
 NAND2_X2 _243_ (.A1(_013_),
    .A2(_000_),
    .ZN(_014_));
 NAND2_X1 _244_ (.A1(CTRL[1]),
    .A2(CTRL[0]),
    .ZN(_015_));
 NOR2_X2 _245_ (.A1(_014_),
    .A2(_015_),
    .ZN(_016_));
 INV_X1 _246_ (.A(_206_),
    .ZN(_017_));
 NAND2_X1 _247_ (.A1(_016_),
    .A2(_017_),
    .ZN(_018_));
 NAND2_X1 _248_ (.A1(_012_),
    .A2(_018_),
    .ZN(_019_));
 NOR2_X1 _249_ (.A1(_009_),
    .A2(_019_),
    .ZN(_020_));
 NOR2_X1 _250_ (.A1(_130_),
    .A2(CTRL[0]),
    .ZN(_021_));
 NOR2_X2 _251_ (.A1(CTRL[2]),
    .A2(CTRL[3]),
    .ZN(_022_));
 NAND2_X2 _252_ (.A1(_021_),
    .A2(_022_),
    .ZN(_023_));
 INV_X1 _253_ (.A(_023_),
    .ZN(_024_));
 NAND2_X1 _254_ (.A1(_024_),
    .A2(_163_),
    .ZN(_025_));
 NOR2_X2 _255_ (.A1(_014_),
    .A2(_132_),
    .ZN(_026_));
 NAND2_X1 _256_ (.A1(_026_),
    .A2(_141_),
    .ZN(_027_));
 NAND2_X1 _257_ (.A1(_025_),
    .A2(_027_),
    .ZN(_028_));
 NOR2_X2 _258_ (.A1(CTRL[1]),
    .A2(CTRL[0]),
    .ZN(_029_));
 NAND2_X1 _259_ (.A1(_029_),
    .A2(_022_),
    .ZN(_030_));
 NOR2_X1 _260_ (.A1(_030_),
    .A2(_145_),
    .ZN(_031_));
 NOR2_X1 _261_ (.A1(_028_),
    .A2(_031_),
    .ZN(_032_));
 NAND2_X2 _262_ (.A1(_013_),
    .A2(CTRL[3]),
    .ZN(_033_));
 INV_X2 _263_ (.A(_033_),
    .ZN(_034_));
 INV_X1 _264_ (.A(_195_),
    .ZN(_035_));
 NAND3_X1 _265_ (.A1(_034_),
    .A2(_029_),
    .A3(_035_),
    .ZN(_036_));
 NOR2_X2 _266_ (.A1(_013_),
    .A2(CTRL[3]),
    .ZN(_037_));
 INV_X1 _267_ (.A(_015_),
    .ZN(_038_));
 NAND3_X1 _268_ (.A1(_037_),
    .A2(_038_),
    .A3(_195_),
    .ZN(_039_));
 NAND2_X1 _269_ (.A1(_036_),
    .A2(_039_),
    .ZN(_040_));
 NOR2_X4 _270_ (.A1(_005_),
    .A2(CTRL[1]),
    .ZN(_041_));
 NAND2_X4 _271_ (.A1(_034_),
    .A2(_041_),
    .ZN(_042_));
 INV_X1 _272_ (.A(_194_),
    .ZN(_043_));
 NOR2_X1 _273_ (.A1(_042_),
    .A2(_043_),
    .ZN(_044_));
 NOR2_X1 _274_ (.A1(_040_),
    .A2(_044_),
    .ZN(_045_));
 NAND3_X1 _275_ (.A1(_020_),
    .A2(_032_),
    .A3(_045_),
    .ZN(Y[2]));
 NAND2_X1 _276_ (.A1(A[0]),
    .A2(B[3]),
    .ZN(_046_));
 INV_X1 _277_ (.A(_046_),
    .ZN(_197_));
 NAND2_X1 _278_ (.A1(B[2]),
    .A2(A[1]),
    .ZN(_151_));
 NAND2_X1 _279_ (.A1(B[0]),
    .A2(A[3]),
    .ZN(_147_));
 NAND2_X1 _280_ (.A1(A[2]),
    .A2(B[1]),
    .ZN(_146_));
 NAND2_X1 _281_ (.A1(_007_),
    .A2(_202_),
    .ZN(_047_));
 INV_X1 _282_ (.A(_180_),
    .ZN(_048_));
 NAND2_X1 _283_ (.A1(_002_),
    .A2(_048_),
    .ZN(_049_));
 NAND2_X1 _284_ (.A1(_047_),
    .A2(_049_),
    .ZN(_050_));
 INV_X1 _285_ (.A(A[3]),
    .ZN(_154_));
 NAND2_X1 _286_ (.A1(_011_),
    .A2(_154_),
    .ZN(_051_));
 INV_X1 _287_ (.A(_202_),
    .ZN(_052_));
 NAND2_X1 _288_ (.A1(_016_),
    .A2(_052_),
    .ZN(_053_));
 NAND2_X1 _289_ (.A1(_051_),
    .A2(_053_),
    .ZN(_054_));
 NOR2_X1 _290_ (.A1(_050_),
    .A2(_054_),
    .ZN(_055_));
 NAND2_X1 _291_ (.A1(_024_),
    .A2(_180_),
    .ZN(_056_));
 NAND2_X1 _292_ (.A1(_026_),
    .A2(_157_),
    .ZN(_057_));
 NAND2_X1 _293_ (.A1(_056_),
    .A2(_057_),
    .ZN(_058_));
 NOR2_X1 _294_ (.A1(_030_),
    .A2(_160_),
    .ZN(_059_));
 NOR2_X1 _295_ (.A1(_058_),
    .A2(_059_),
    .ZN(_060_));
 INV_X1 _296_ (.A(_199_),
    .ZN(_061_));
 NAND3_X1 _297_ (.A1(_034_),
    .A2(_029_),
    .A3(_061_),
    .ZN(_062_));
 NAND3_X1 _298_ (.A1(_037_),
    .A2(_038_),
    .A3(_199_),
    .ZN(_063_));
 NAND2_X1 _299_ (.A1(_062_),
    .A2(_063_),
    .ZN(_064_));
 INV_X1 _300_ (.A(_198_),
    .ZN(_065_));
 NOR2_X1 _301_ (.A1(_042_),
    .A2(_065_),
    .ZN(_066_));
 NOR2_X1 _302_ (.A1(_064_),
    .A2(_066_),
    .ZN(_067_));
 NAND3_X1 _303_ (.A1(_055_),
    .A2(_060_),
    .A3(_067_),
    .ZN(Y[3]));
 NAND2_X1 _304_ (.A1(B[3]),
    .A2(A[1]),
    .ZN(_068_));
 INV_X1 _305_ (.A(_068_),
    .ZN(_166_));
 NAND2_X1 _306_ (.A1(A[3]),
    .A2(B[1]),
    .ZN(_069_));
 INV_X1 _307_ (.A(_069_),
    .ZN(_200_));
 OR2_X1 _308_ (.A1(_030_),
    .A2(_159_),
    .ZN(_070_));
 NAND2_X1 _309_ (.A1(_026_),
    .A2(_156_),
    .ZN(_071_));
 NAND3_X1 _310_ (.A1(_034_),
    .A2(_041_),
    .A3(_169_),
    .ZN(_072_));
 NAND3_X1 _311_ (.A1(_070_),
    .A2(_071_),
    .A3(_072_),
    .ZN(Y[4]));
 NAND2_X1 _312_ (.A1(A[2]),
    .A2(B[3]),
    .ZN(_175_));
 NAND2_X1 _313_ (.A1(B[2]),
    .A2(A[3]),
    .ZN(_073_));
 INV_X1 _314_ (.A(_073_),
    .ZN(_170_));
 NOR2_X1 _315_ (.A1(_042_),
    .A2(_178_),
    .ZN(Y[5]));
 INV_X1 _316_ (.A(_182_),
    .ZN(_074_));
 NOR2_X1 _317_ (.A1(_042_),
    .A2(_074_),
    .ZN(Y[6]));
 INV_X1 _318_ (.A(_181_),
    .ZN(_075_));
 NOR2_X1 _319_ (.A1(_042_),
    .A2(_075_),
    .ZN(Y[7]));
 NOR2_X1 _320_ (.A1(_033_),
    .A2(_006_),
    .ZN(_076_));
 NOR2_X1 _321_ (.A1(_195_),
    .A2(_199_),
    .ZN(_077_));
 NOR2_X1 _322_ (.A1(_213_),
    .A2(_222_),
    .ZN(_078_));
 NAND2_X1 _323_ (.A1(_077_),
    .A2(_078_),
    .ZN(_079_));
 NAND2_X1 _324_ (.A1(_076_),
    .A2(_079_),
    .ZN(_080_));
 AOI21_X1 _325_ (.A(_203_),
    .B1(_061_),
    .B2(_207_),
    .ZN(_081_));
 NAND2_X1 _326_ (.A1(_077_),
    .A2(_139_),
    .ZN(_082_));
 NAND2_X1 _327_ (.A1(_081_),
    .A2(_082_),
    .ZN(_083_));
 NOR2_X1 _328_ (.A1(_080_),
    .A2(_083_),
    .ZN(_084_));
 INV_X1 _329_ (.A(_186_),
    .ZN(_085_));
 AOI21_X1 _330_ (.A(_085_),
    .B1(_042_),
    .B2(_023_),
    .ZN(_086_));
 NOR2_X1 _331_ (.A1(_084_),
    .A2(_086_),
    .ZN(_087_));
 NAND2_X1 _332_ (.A1(_002_),
    .A2(_085_),
    .ZN(_088_));
 INV_X1 _333_ (.A(_212_),
    .ZN(_089_));
 NAND2_X1 _334_ (.A1(_016_),
    .A2(_089_),
    .ZN(_090_));
 NAND2_X1 _335_ (.A1(_088_),
    .A2(_090_),
    .ZN(_091_));
 INV_X1 _336_ (.A(_213_),
    .ZN(_092_));
 NAND2_X1 _337_ (.A1(_037_),
    .A2(_038_),
    .ZN(_093_));
 NAND2_X1 _338_ (.A1(_022_),
    .A2(_130_),
    .ZN(_094_));
 AOI21_X1 _339_ (.A(_092_),
    .B1(_093_),
    .B2(_094_),
    .ZN(_095_));
 NOR2_X1 _340_ (.A1(_091_),
    .A2(_095_),
    .ZN(_096_));
 INV_X1 _341_ (.A(A[0]),
    .ZN(_210_));
 NAND2_X1 _342_ (.A1(_011_),
    .A2(_210_),
    .ZN(_097_));
 NAND2_X1 _343_ (.A1(_007_),
    .A2(_212_),
    .ZN(_098_));
 NAND2_X1 _344_ (.A1(_097_),
    .A2(_098_),
    .ZN(_099_));
 NOR3_X1 _345_ (.A1(_010_),
    .A2(_033_),
    .A3(_213_),
    .ZN(_100_));
 NOR2_X1 _346_ (.A1(_099_),
    .A2(_100_),
    .ZN(_101_));
 NAND3_X1 _347_ (.A1(_087_),
    .A2(_096_),
    .A3(_101_),
    .ZN(Y[0]));
 NAND2_X1 _348_ (.A1(B[0]),
    .A2(A[1]),
    .ZN(_102_));
 INV_X1 _349_ (.A(_102_),
    .ZN(_217_));
 INV_X1 _350_ (.A(_189_),
    .ZN(_135_));
 INV_X1 _351_ (.A(_083_),
    .ZN(_103_));
 NOR2_X1 _352_ (.A1(_103_),
    .A2(_080_),
    .ZN(_104_));
 NAND2_X1 _353_ (.A1(_041_),
    .A2(_037_),
    .ZN(_105_));
 NAND2_X1 _354_ (.A1(_105_),
    .A2(_135_),
    .ZN(_106_));
 NAND2_X1 _355_ (.A1(_023_),
    .A2(_189_),
    .ZN(_107_));
 NAND2_X1 _356_ (.A1(_106_),
    .A2(_107_),
    .ZN(_108_));
 INV_X1 _357_ (.A(_108_),
    .ZN(_109_));
 NOR2_X1 _358_ (.A1(_104_),
    .A2(_109_),
    .ZN(_110_));
 INV_X1 _359_ (.A(_221_),
    .ZN(_111_));
 NAND2_X1 _360_ (.A1(_016_),
    .A2(_111_),
    .ZN(_112_));
 NAND3_X1 _361_ (.A1(_037_),
    .A2(_038_),
    .A3(_222_),
    .ZN(_113_));
 NAND2_X1 _362_ (.A1(_112_),
    .A2(_113_),
    .ZN(_114_));
 NAND3_X1 _363_ (.A1(_034_),
    .A2(_041_),
    .A3(_219_),
    .ZN(_115_));
 INV_X1 _364_ (.A(_222_),
    .ZN(_116_));
 NAND3_X1 _365_ (.A1(_034_),
    .A2(_029_),
    .A3(_116_),
    .ZN(_117_));
 NAND2_X1 _366_ (.A1(_115_),
    .A2(_117_),
    .ZN(_118_));
 NOR2_X1 _367_ (.A1(_114_),
    .A2(_118_),
    .ZN(_119_));
 INV_X1 _368_ (.A(A[1]),
    .ZN(_220_));
 NAND2_X1 _369_ (.A1(_011_),
    .A2(_220_),
    .ZN(_120_));
 NAND2_X1 _370_ (.A1(_007_),
    .A2(_221_),
    .ZN(_121_));
 NAND2_X1 _371_ (.A1(_120_),
    .A2(_121_),
    .ZN(_122_));
 NAND3_X1 _372_ (.A1(_029_),
    .A2(_022_),
    .A3(_188_),
    .ZN(_123_));
 NAND3_X1 _373_ (.A1(_041_),
    .A2(_022_),
    .A3(_185_),
    .ZN(_124_));
 NAND2_X1 _374_ (.A1(_123_),
    .A2(_124_),
    .ZN(_125_));
 NOR2_X1 _375_ (.A1(_122_),
    .A2(_125_),
    .ZN(_126_));
 NAND3_X1 _376_ (.A1(_110_),
    .A2(_119_),
    .A3(_126_),
    .ZN(Y[1]));
 NAND2_X1 _377_ (.A1(B[0]),
    .A2(A[2]),
    .ZN(_133_));
 INV_X1 _378_ (.A(_173_),
    .ZN(_176_));
 INV_X1 _379_ (.A(_140_),
    .ZN(_155_));
 INV_X1 _380_ (.A(_168_),
    .ZN(_174_));
 INV_X1 _381_ (.A(_187_),
    .ZN(_143_));
 NAND2_X1 _382_ (.A1(B[2]),
    .A2(A[0]),
    .ZN(_127_));
 INV_X1 _383_ (.A(_127_),
    .ZN(_191_));
 INV_X1 _384_ (.A(_153_),
    .ZN(_196_));
 INV_X1 _385_ (.A(_177_),
    .ZN(_179_));
 INV_X1 _386_ (.A(_214_),
    .ZN(_184_));
 INV_X1 _387_ (.A(_137_),
    .ZN(_192_));
 INV_X1 _388_ (.A(_148_),
    .ZN(_201_));
 INV_X1 _389_ (.A(_152_),
    .ZN(_162_));
 INV_X1 _390_ (.A(B[3]),
    .ZN(_158_));
 INV_X1 _391_ (.A(B[2]),
    .ZN(_138_));
 INV_X1 _392_ (.A(B[0]),
    .ZN(_211_));
 NAND2_X1 _393_ (.A1(A[0]),
    .A2(B[1]),
    .ZN(_128_));
 INV_X1 _394_ (.A(_128_),
    .ZN(_218_));
 INV_X1 _395_ (.A(B[1]),
    .ZN(_183_));
 INV_X1 _396_ (.A(_193_),
    .ZN(_150_));
 INV_X1 _397_ (.A(_190_),
    .ZN(_134_));
 FA_X1 _398_ (.A(_133_),
    .B(_134_),
    .CI(_135_),
    .CO(_136_),
    .S(_137_));
 FA_X1 _399_ (.A(A[2]),
    .B(_138_),
    .CI(_139_),
    .CO(_140_),
    .S(_141_));
 FA_X1 _400_ (.A(_142_),
    .B(_138_),
    .CI(_143_),
    .CO(_144_),
    .S(_145_));
 FA_X1 _401_ (.A(_136_),
    .B(_146_),
    .CI(_147_),
    .CO(_148_),
    .S(_149_));
 FA_X1 _402_ (.A(_150_),
    .B(_151_),
    .CI(_149_),
    .CO(_152_),
    .S(_153_));
 FA_X1 _403_ (.A(_154_),
    .B(B[3]),
    .CI(_155_),
    .CO(_156_),
    .S(_157_));
 FA_X1 _404_ (.A(_154_),
    .B(_158_),
    .CI(_144_),
    .CO(_159_),
    .S(_160_));
 FA_X1 _405_ (.A(_161_),
    .B(_162_),
    .CI(_163_),
    .CO(_164_),
    .S(_165_));
 FA_X1 _406_ (.A(_166_),
    .B(_165_),
    .CI(_167_),
    .CO(_168_),
    .S(_169_));
 FA_X1 _407_ (.A(_170_),
    .B(_171_),
    .CI(_164_),
    .CO(_172_),
    .S(_173_));
 FA_X1 _408_ (.A(_174_),
    .B(_175_),
    .CI(_176_),
    .CO(_177_),
    .S(_178_));
 FA_X1 _409_ (.A(_179_),
    .B(_180_),
    .CI(_172_),
    .CO(_181_),
    .S(_182_));
 FA_X1 _410_ (.A(A[1]),
    .B(_183_),
    .CI(_184_),
    .CO(_139_),
    .S(_185_));
 FA_X1 _411_ (.A(A[1]),
    .B(B[1]),
    .CI(_186_),
    .CO(_187_),
    .S(_188_));
 HA_X1 _412_ (.A(_191_),
    .B(_192_),
    .CO(_193_),
    .S(_194_));
 HA_X1 _413_ (.A(_196_),
    .B(_197_),
    .CO(_167_),
    .S(_198_));
 HA_X1 _414_ (.A(_200_),
    .B(_201_),
    .CO(_171_),
    .S(_161_));
 HA_X1 _415_ (.A(_154_),
    .B(_158_),
    .CO(_202_),
    .S(_199_));
 HA_X1 _416_ (.A(A[3]),
    .B(_158_),
    .CO(_203_),
    .S(_204_));
 HA_X1 _417_ (.A(A[3]),
    .B(B[3]),
    .CO(_180_),
    .S(_205_));
 HA_X1 _418_ (.A(_142_),
    .B(_138_),
    .CO(_206_),
    .S(_195_));
 HA_X1 _419_ (.A(A[2]),
    .B(_138_),
    .CO(_207_),
    .S(_208_));
 HA_X1 _420_ (.A(A[2]),
    .B(B[2]),
    .CO(_163_),
    .S(_209_));
 HA_X1 _421_ (.A(_210_),
    .B(_211_),
    .CO(_212_),
    .S(_213_));
 HA_X1 _422_ (.A(_210_),
    .B(B[0]),
    .CO(_214_),
    .S(_215_));
 HA_X1 _423_ (.A(A[0]),
    .B(B[0]),
    .CO(_186_),
    .S(_216_));
 HA_X1 _424_ (.A(_217_),
    .B(_218_),
    .CO(_190_),
    .S(_219_));
 HA_X1 _425_ (.A(_220_),
    .B(_183_),
    .CO(_221_),
    .S(_222_));
 HA_X1 _426_ (.A(A[1]),
    .B(B[1]),
    .CO(_189_),
    .S(_223_));
endmodule
